XlxV64EB    1ad5     9e0�͒�6fxf�'n�mẅ́�i�PWa�[��P�HЉ�V��7�G��fF��~����w�q�nk��P�q?��aPb!�:�#�!�y	�C~K�t�K��\��s��J���J��H�yW� k�GȪ,���
9xJ�@��<v,~�U�,�;�+W�t:��� n�
n� ���\��%��"����D���d+;��U�%��zf�Z�`H;2��D�����0���e�׸� A`�H69�d��cΈ���$��t��' �9)�=E�qP��2�l�01R�G:b�|@������$iQ�j���6�=q����r�؛W���]c������i���g�j?k�A�1l;q?h�W=XO��L,�0��ѣ�8"�����a���U<���?|u3����xz~����+��V�����jM�U��ޞ$:�1OA�l����G���E	�>ةb$ؒ����hÈ�F�l�l�$<%z?�w���O��v��2���?UE���w�,h��XC�:�>�THHAOS�į�A��ZCt}B�Mz+V5_��l�:�<5�Z�����|7~k�����٧�G8\H�9>ԍ��H!���Z��D7,�J�Uv�����y%z�^j:/�en[]f�f��Fe��ֹ��Ш'���Yv�[�@-=���#FxK����H��`47����b��oY���ʂ�\�	�AW�J��B��K2/�r�e$�@��m�l#��Jz3 !��k��Sz���J?���B\�Zt�~}�q�"�2�^#��A� ���?TN�'\�I�iI���po?y�����#��oXE'3��-��k\�̃���ۮ����D�╕3�q�(F�@W<e�eu��	�\���r�.~_��ɭY��2�*��ў�w$�ň��j	����"�O��=6�^["}�����cW�.?@_��4�f6[�����*Y8(�����.��A���s}s<!�;nU{u�!�V@l��ր�}]��Зo�_C[�c)�k�/N+&8z��YΌ�{L	�+7ӯ��妻{��j'�v�4Y��(�f� ��e�"0�F��]?�g1�d�ͳ���ċ)��G��a�7����p�
�"LK���dT�'b�Ϫ����>Q��ƥ��him��Cn�Z��bbޓ:uf��]B:=s��@�cG^���Л�r��b��W`L	t���˗�֤�b��i��0o���X_nc{G�8�72]�?'�t��!���k;y� V\��Gn0sJ;]a��޸>:?>��rA�"�u�**,��:h�� ��3%���F*��0�`n�j��u�ez}LQL��kAʕkC\CX�~1α�2)+2|K��?��>���Le(ȧ��!����e�1�����k�巔��zu�ϣ+: 7�"c�:��Q�)Em˖Bbq�{��7�(�JO��/ʨrM���6$���|�~��4�녊-�!����ΝGcR�/�@[�z��^�_�P\`&�8 �'T�7<2F��_Zsº�8�g�f��.�O�������:S����;jI#?�8^�em��a�0x%ssr�XC¾��*��)� ��?�q����Y��=5�|�<�ˏ�u�u�Ȯ���&eV�l��wc��h
NEBqV��#�V~�;�gi/���A8zᄕE��{[��sG�EZR`�{؆[������0?��%פ����>daq{��(�^�ξ[����s���O^b&��"��T�^��^��{�0��u�kP�����'-���Kd�V�x�m7
^�>���� [[�N�(�4f�t����5�?w�w�	D8H�n`�O�1 !��WǂLfՈzl�!�������׺�>��uO���Aߴ�4�:l�b]��J@�7g�?�#S$('���	B���@~�\�i�:�AȦ�zá��N:R;=Ak�ZK·EL���FB�%!������C��OW4s�J�+3ɚ?�>-������M)Y�ͽU�/���Y�y�ڸ~q=�ݤ �6��n�;-r�����)�{��N���g�2vp�PQ�%�B\�m����!,UN ���/�-%\��|��r�@�n���;���[34�ߊ�=��aol��2	��%��i[�OR`"/]^�&NX�#me	�ޯ�
���+lg[��ĺ�<�>=Bn�yVȈ��2u�%j��a�Z���׆�6A�5�.V{���ƛ������37jr�hPR��r�bX6�mG�D.��6��}c�����H�GLE	�^�-���4�Ix������b���UJP�u=�O�E�*۵XW�Td��H?�sN�:���Ǉ�/C�`���s��rV����c֝0���-�����|o����K�����L�����>e�y�72#�,�M�B�زk�����gPR;�|j{���K{AM�c���if@��j�cF�B]��N��:�6���6����5sV4�X���ʇi�N9hn�g��^�yz��0�.RJƴ�