XlxV64EB    823a    1470�on]���fjL_�&�jE�p�륈v�o�qX�M�OSx����y/���ɫ
��&��G\����{6��4�����N'�Y�2�4uM��{̾s{���4/����� -�����o���@�3R�ϕ�p��N՚:$�e�-E&��|�:=DB��E��n4��J�!�ZqcsW)չ�<v�}Ċ-&C�F��䙷l�jl�N�V��I�7�Yԟ��"�6|���볩0�S抶�k/�D<j�*y������j���~��`��	r̞��m���Qf�{^��/��:�y�` r�����٤QE;�K����Ű��uO,��fᷥ@zX�^�S}�eՇ���B�z�N5U$�L�#�K{����OG���W���e3�8iO�s��6R���JF3�mc��q8z8�6�d����9��0]ֲ�gp��^�]<qn*{�اʋ�Bvd��<��}:�dԚ��L#5�*D{َ[�&� ]H�u��1�F��V������p�%��ڍ'���4���R�j8g��*zB�rY5~�����Сz�0�\���LH5���{� 왰���㚝\k�.o�p
�,8/(�{����7߬��j��4����=`�h�mLK�:�p��v��N�V��e�
m��,5��9��W�C� �I�^x_3I���I�z���Fy��*�2�H���Ƕ���&�! 9")�i��WL����ƀ�h���?��)���7�#�y�ֳ�b���pcN��
����U���6�{�Ы~�
Ⱥi1��I�.�	��/�Aϛ/Ŋ�؂�Y0��H�?���t-tq��9��b�.l�U��9Q$�'���oS^nzR攅b��lˎh�>��7��~�C�rd�7��n:�&��,5�W������
�2�1��bщ��EҖۿ��ۗ��%�-UC�G>l�Y�ߢi�o�[f#��L�Y%ް	��OI\(��G�sTdCl�L�9�G��ů�{�L n`-Y�ׯ�_��t�k*�_�!&)����6M�	%؃�����}���vJ����i�p�ݜ���r��5E}#���`ފ6B���F�2�8:3%W{<�-����аB-i՟����b�bGK�`��3X����բR��,!����3f���*�|N� �Q8S	���O��E�����������E����`�x�d�v
=���x�r���B>>|��6�mR�G�ޟ)�H�sH!��$ťQ��6�~��<�M��	�[�q� ��h���P-�~p���I��T-��BvO��;��˸h+Y��u(h'��N-��v/��<�� �r:�$�~8��	�XB%D�w�\����7��x��Vm�@K�(���=�����ޮ_�{{�4��d�屇�}��\_���/����	yő���K>#�k嫦�����Ց倡mx��2�or��T��r��ʱ�_[b�Dȋ�}Fċ�y��@�Ǖ2���)|KWV��Dx�K�op�2ޏL.�?�6 �'���5��[x����ʎy���o
���g��S�g�Hlw%�;!f\��I�SS��y$3�߾�|�I҈Ec��2M���I�i����I(��)z����j���|4�D8,=|��8%���-m���ǔ�O�9Q'!<f���5U�IH��-q#�!�TuN���V�Q6c���k��a�yۮd�[�k8��,�C����sʪ�/���������s��/5٢����L���XLІ��U�.�fE����2�Ǣ��uْU���4fl��p�^�b�11���3�y���}ف�w
��
%��/�w��a��+��3V��:�k �p��QH'�3��I�r'"�{��~j-Yq�b�92��:��� k������D�Y��j��_c�4���mZy�	�1�+��pi1G�0�.�#DS������M���������$惽7�`	�\��μ��+�<5��h䧇�`QV��~@��Iȣpa/p��y?��	�ה��~;�Hڗ���Q����y,�\m^��o�r�n�3��М�I�h��@�Ϡ���kd�Ⱦ�e�55,���w��ǟyO�bx�[�1l6IERqc�VZ����2E��=q�,�Z O!0���Z������Q�{�2�0X�P��(ى��h�dLB5d��JH�_�1�nף�N8]Fhջ��X�31'SW���p��gC@��/m���;W[���{��[�(����h��$��x2	O��,��Q�J%���z��'�ӛz���x�5�C�*4�6��'�Q\u�%�ze�4Tub��^��˼2�>_a[Ž6�t���ELal�!Ͻ~�v�	B.u�1%�2;�GL;��9��<.)a�h)A�H*$�l-� �$J&����L}�� 0NrF�1�*��|�цhm�v�I�q�{Q�B���z���.}~�$�+��)(@��Ƃc��c�kڶ���ۺ�����@���a�`9�1
���0���q�9�-��14�`ѻ];��7�@H�����P5��8��^������5���B�ń��oX�R��\�Q�889o65[y<�"U�l�Pm9"/tT�A
���FhI��e���-�������'}C<�6��W���K�k89�/)#_�]ݨBǊv􇜥ik-��SeqtK����)K=qbw�-�d,�-.�PE�Xa��:�XC5oX���W��UR�16�3��R���{�	���)\-�O	��k��b`������(uϘQ�����lg�Z���Ɖ��?x�"bi���;?������'7H�QJ8�C����n���Q^hd��d{i옎:q<�i.�2
k݂�D��\ ʚ��ӫ�����oN�}3��.1�<�N��>�:�(�t	>�,�(�[�6购�̇�ͩ�D�C\X���I��u������.�2��$�~��!9����T�ZM�ڋ��KT�,M�悯x�w����"���N}[�~��Y���ɨ:���&+b��R��fZ�@:�U�_�
��f1�k���C��X%� nA��Cl��sդ��s�@�/|W�!`sD�m4��2�1�T�*!���V�Qr~ܑK��k������I��D��l�����t��9~*�+�Hb�{�LZ�+�d��J�-,��If��ȷ�=RZ���,4���O�Ԟ�������#F��Zp�v#�ܮ����?�{�o���$@����y���ZҚ�h��["C�
7C�U�v��NR�Vv��
8`F�����`�������h`H�tG���lBtF2ƼBPe��2��$J�D	�00�V�n��>�zX�N�R�Ї<WR�7��c:t�}�"&�ھ��a�#�9�ˇ���V~��Z�]�u4k g�+��$�i-\D#���),�nS٭
S}L����;��^\�O-��`�����J76��.c�g�(1�gu9/7)�6o��B��1!�Ju�峓Х���l�V��.�.�"�y4�q�X���"%8�Ŋ�(�4 AAY1���\Å~"ur�S�4�Z���{SAb-nNAO�2�	R#?jÖ �徱����ieZwz�j�u묫v�'7���u���J���o� �#Ui<��K���D��asc�X2�q�w3D<��}8�@�����`�1P�F�{���ۆ�_L�W�����Gs�<�	}��jf)�@j�n ��A@�勌����o��}9T�W�f42v�N�ܢ-q���G��hD#	ߗZ"P��^X=O�HM���Q��e��:W�8�B�Ͻ����{��(���gp�_��d���o.�yC�6T1Q���#�Z���]�j��Z��F]>����JG�B	��<�|�#0�ܹn���HR?f�[*�o�/��V�F
�n�<����%Kg�]�I�	�ʤ�:|�����i�X�����l�"a,�m�����`��|'��慥k�;O��ɷ�f�R=id��ؘ�;w_"� E�ʻ|�G�l�x�Ja³�{-�W``�^讥��Q^�W��c�f��ޅՎ��_���Mi��\�?�&1>(�*�B��K���S6���JD�a�x��R��(g��)�sU 4��΂X1�lo�\I�Z�BK�w��e<���Y���u���b�?]������Ny���Ĭ�)�mLc����8y;���9[IʾJ�G���8t�c-��k
��Vj*�Z��T@ �?�����ҏ����8Ӟ�9�,��uJ	�b�@����Q�_�.m�v#�2��]pd�٣I��%4�E��8��	�"�U�WQ��c�������[�y��z����G̐��i�ؗM��(��$�%1��%�W��'���xSg�T_� OYF��"Ȉu�'.+2x�OWU�#���yH�L`���`�	�B�����?���u>��3/"�����H��
��W�|5���0��*�/$�w�k��߮�a8{牢U�� C�ET]@�4?�9Pr��*s?.�M�O�.��������Ի<�B��Z.�9�w�FJ5j�{����Z�ΪB��Uu^�*,�4�K���Y���:�3D(F�hK�i���)J�w�YC ȟ���	U�~��#����e8��sr�4̈��'���ZV��Jh9�嫖*�j1��5����[�mo2<+��C�ηVM��i0p��j�A�G!wX�� k.�Ba�oa$���>��!8�W�2�h���/k��se��w�/?��,O��%j�_���ғ4����{!�<*��C�S@�Ő�:'�<+y��؁K@���o��(A�臗̥a��NX�������pM6�Њ7#�l!���j�47�Ժ��d0�C5(�fM1���]q8~�ۊ��ۦ[b��[��	�0���c���FH���7`�U-	H5n�C�I�r�)�\��]�ه�-�ih�|B7w�˗�[�v�ZSAH�'��=�.~xZ7���_Ia�]͖h\2Yu�L;��م�\-<��ٴc�iҲYv>��v�eP:^A�*y峺Ƭ>���Į s��	��Ry�w<]N�t����]�q��T���}2��3Q#/� ���"9�'�7����cK�I��v��M{V�����5�V�,�o;RZ=�:t��p��s�`�&ȊSƘH���|��|Qq�������(u7�*���=��P�R�oR=�����u����