XlxV64EB    1f73     9d0
�)v#�5ŸP/ ��~�v>#�F�Ƶ���D"Dw������JqX
i�`;+�&���&�3�ͺr�z�kb�����ũL����~��iV�@"���kz��8�yy��i���P��u�Q��6����)�T���{��Λ�tE� y���ҡ˃H��Q� ]���־�i�jJC����;�Dֲ��G=<�:Z�S�jl߿`k�L$*�d	_�	5Zb �<h�bwD��Oڲ6q7e9.F�j�����8��2/�킗>h6#��
��j�ZR�����u�L|��w��}T�S�֢��6Α4�I��*�<�d ������w6|��ٖ+�i3WRi�`E��dF�~⾐��R��~0*]t�'���v��&(j�C} �%X��V�����H��O���h+�SW��#%���{���H�Z�;�;C�{��>�z]_�}.FEQ�'���uʏB��X#���Q0F����%G�5A�7-������!�fzv~�P��T�F�.�>Wu.Q��+��6DE*�����G�MS՟r�-�v��4l�t7օ�D�L���G��!֛��\��apm��Cי4�'�(yQ���9����7��<n)�0+��9 Y�6�67s��5�#U4������ND�I��;�U<{�U�#�	a@��DpG�f�׻&w���a��Q�`�����9E��7P}2�e��X%{�1����%]��[�_p�D�y���"˽k�o4gisIΞ�}hDר�Z��\GF��ǟ֚�,��k<'�;A�����I��N���D%��U�D%8a��4��"V��5)f$3��Bؿ_$�d��E��l��3�F-^
�쯰�sI��w:hx�oX83�� �*���t���y��C'��G��D���K�#�3��Y��RqC�{2����M���7�J%g���ػҩ��?�_M�KL٪�����������#D])�R'�������X�{��@�Ǐ����o�p��{	�rq-���1~��73K^�W׋��e���K�E��
������Gؘ��2�%��"��k����Ssk�e����e+�c��r�eOLd��ҍ���Q�����V�"�O�$�N��dzUr�cוbr��"�]����������[$�0��]�<֓_�ɋ�.ͼsfV�Y
�h=����5�	��[:����O�t�"����9��0����Uځ����f�5�!X�gQP8�%���nA�'[Y������p�Nϧ��Š�bm����}m*r�� ̶��L����]�W�Y���^H��S����S�����\�@����ԧ�v�(3-����w��)�f��  .B#��4���萬0=:	�s���m�hJt`�\��B2���<��
S���[�ؽK@f��/l7�׭�����4iӖyf�DL����g¹������D�yW��D�`j��ˢPqh����y7������Ӡ�g��[M>�|���]B�_Ia����i�[I>e�8��=�B�9�d��؅�X#,}U"6�PP�>u	����!E�H���ct͐]���:���G�AP=����H�Թ��ro����*��~H�����w�7��6�<��y��Kl�q�QȞwB�Ȳw���v�6�p�R��Ի���N�6&��+G��P�V��-9�4M��!+���L1H�^Uߖ565��6�U�;n(�1�� ���yW��s&1'AŽk�+�[�&���#A� )p�)k֊��^���:&[�m�CK�dL�"�<%2	���� ��W�17�4���>k��� y����#�|��A$x����N����:�ZJO������؈�k���b�U�*#M��x�z?c�][��� jl�(<��od$F�Āh�M��O>I��c�� 	^�G�H9�_���֒\�qV �����{]Su�Ϟ��B3�B`[���rѡ��ugE��(Px\�Gw]ɍ6ᭈP�"�nR�h�.������ەa��c�PiV]��e������X��~�Q�&I%�D�a��T�V��L���0�.��"_��MO�OC���:�2��`U���!�xn��ID�c�a;a�R#�[��w��<���-��%��e�}%{����)���/-�F�f�dێytт������P`l>�S,�7+�����ݳ1Z���z�W\�W��Y|+"��,��oFh��}L�Xk��w�q�����HA�'&*�`�R��%��=�u��:
�hfc��I���j�i�ɾ�Ct�\������0��m�;����s�t5�c�_�� Ւ����q�OI[�oϤ��Mgx0ڨ|�%.�*'\�S��o�m�`Ӥw�^쿉���'IC�4�*�ZF㗨D҄Q��-��c�ཞ�n�_:�+���>�6���Y�$���脠�$�q�HF��lV[�e�&؀Kkz��-�R��|�7�[�DJ&8��#)����G�|n6۹?��e�;���L�b8�z�b��Կ�