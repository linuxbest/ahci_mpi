XlxV64EB    4910    1170T=BG�;Y��X5*����m*\H�w�ߋ-	��<���3. g�i6����w�l�O�o
�C�m���|	����W��ە~P�/����N%𔿗���[��D�)!Y�6**AQ��U�TN��i��"�S���Ǘ���D�A�{�X�r,�G�]p" ��A�U���4UhYs�ߵ���O�¤�*l���Bi��֭B��;_���	e��D:�O`)
ࢄ�į�WB��n6ծ,�2�'Mv5mC^�����.ܝ���<o£Ѡ��	�a�ѫWv�I�V�y�}�=�?�gW�t^MVf����J�-b�bӼ!N��� V��:�F4besu�����_vL|��=�V�u�+��ZJ#�zO!"z
���9-�]����0+�R��ş��O@�46�N B/5e�ɺ�L�P�k^������5����R+:p��຃ю6�87���v�C��^,N���A9o��w��~�p�1<$h����U��6�����n�c�����j|��i��A���Q�'PHs-����j,�JH�������{r���n��+1�uo��"g7��V ���&l��'�ZXM�����v�H魺&����
�XQ�e��'׉�W��,����{��(ek3R�=�g{# ��a�6�K=�>H�Z�l��)�b�^%�J"���"�ܰIty3-��?�Is�ڏ��0[\Lr��Τ6 >X�m/cm���,o�f�`L�ؒj�1?���� ՠ�k�X��F��Be.d�����>p(Y_<7�z�����:�z�l�b�U���,`�he���S�q����)�e�F��WO���
b	g�Rf\m�ю�?��ރ��!J�V�'�p(X���S���f�QΘ�42Iݙ�>VƳf�c����+��>��e��>;M����3k��M�	�J!�{��w��/��r�[�c-��
�B��{QY@6��HHK?�hd>r >�\�i����*"֪^�!��J+:٘�9	�U��΍F�I��i]g�h5U5N�����#��s�v�����C(B ���]���m�-�$r�l�d�Xn�n�-�O��,mFR���`�v@�'C��ct���L��q�C�m�.]x��ݼ��m8�#A�_��<َ���$��H����@��:�e�W�,R���x�*���{��ws��Yxw1
0�}Z��tY�����~�7�gj4��G_+�(0���&�Ϊ�XzP8��+�\#���2�z��������V��.�s��%ZJ�(����e9Қ���IhWw=ڏ���<���1?�'ϧ�S����d�(��F��e̘d�"`n+rE(P&�zv����Xc0�+'!�����h16�|�x��2�/�q�`����J�x�>���c_�41��2��-V���g�lN`��@h%����7��b�䮒ȆH��޸�bQtb��#/��P�$��0��5[�l4�*#�0�
�=��.��|�y��>�P�Y�@Bxz����z?z~��
iQ��4�j9En��b��/#�쿵������-�<��c����߅Y�s:���F�Lt��&d�8��<��;�`�Q�u�X�dQ"�v�&+&dh��d��Z�x���検>�lu)��l��a	!�QU��ʶ�� �볱��&W�GG��v^�-���u%�.�ŧSS�R�'��	�,��r��N\�_��]�!-}G���h?��͍�<�$�8��t*t���ey�
�
���ǖ�9S����U�iJv��ߟ�� �a��,�ܮF,}�e��T��-P�_��j���[����TbMdDE�t�������#S������&����?c�6 �4KF1Z��$~:���ָ�*�d�2U�V���kW��TA�9�227�6�·�A�ĺ��:=�\869/��kݮ��b�����Hv]YE"{���s�zݧ	��з�5�D�PF^yz�v���0����c��K�L�vQ�"Sn3�I��T0m���
�`����W���N��H]7�g �;���
s�8u��6�������FT��	ʆ��)n�T��ե�f��������[5C��ټ�0��:ڔ�j]�N�SF�l�:`�d|}�}���o��`�`]1�-���M�e��Y���?��4�)����I=Z:F�QH|%�aU:M,=\�U�)O����ʏ����EZ�[��eQ�M��#�>��Ug_YI0�Ϥ�6��w	��x���YY���5@D��B:���.4��T����~��pm�ZYM��%]��w6	�;�ho�r�&LU^ˏ_�Pl�^{}�+ۋ@�Tj8_�	�&�`���ؾ��i���T�w�jz�i��/.��Y��-f�N_,�����Sm�{Gs� ��=����l������]m3�cH�
��ܦi��>��wCTCN��aڍ:mk8�J�ɺ�.Ug��YD{��n$fx�.��ܓ����P���]k4$��L��k�-�;B�0��膰Ո�<���J�^��`C#������q&|'������M�y/+��#�b:�oh|h�Yˈ��'��}�-��W�'��C����=�V���I�\���7勛�J�V��׫�>��5���4����1/Ii?r�,��$�ۦ�:7�M�����+��}I`��Mظ쭁->d~�|��t�Mf?���eq�4�f`�W�#%[=�2q�ɱӥ;�!k^����y�t��#��I|4�M/\є�P=7��e����D% ��SG`�j�Ϗ��8�~�ڝ��u������uLґ*��?V�9�E���e�.�5;'�G�_�hՖ"�23�H\�*,S�#��gK�@tI�t��H6`���S��YPz#koo������PEӱ��$ޛ�.�1�y���6��_��z�0��2&P|»3��τ�`��c%�&��?єT(M	������Dv3��u�~��$��
�����e�vO\ul�2&#��B��>���F,J YS7�T���g�����I�8��V�?h����c��5��T4�W2�-ȡZ-�p�i����O�q�׺؟�!RoYA�G���⾔�e@�>�I����Z�A0ۜcW` �a�r����� ��L�E�]�ኒ���RȥBZp,�~�����d�]:�9^^˫�� �J�!-.�xIًd�f�"���Yx&���0�i� 5*?��z��?������Y���/����J>Z9�J&oXӞ,L�\���/�t�l"���`���_� ҥ���MV�B�єKH��
��t�?,��Y�!r�u�~b�i�Ui�9��bZ�H�c
�z�!k	
]2hȵ�}5��7(��[erd��7m�'*0C��u�^�_$��`�B�����!�?��)�b̆��q�&��$�j�q��1�b^'A�e�{I�J��2�\/�h��}�͛:.JS�X�][�T������4�*^���UOx�_~+��SBoa�Y1�8��R%K3䮖���M������N�'�&5�4E4=�FA(?t3��sv1���c$`Onq��TYȯE��pȻ_���|/fg��J`�3�	�{r~�R(י�8���Z~�
	��앷.��s(�X��Jӥ=��n5����uL(�-�@^ u���2Q�S��s���4ŰMdާGH1]��H����-�e���wmX��rq����2��w����'�PӢ��5�c8����u��I����]��*m!��oMI�({ӽ�'E��(���#w���©�Cn�,��C��������M�q�;��j�Pg����4�mY�QPM�t9$ʹ���9������}�80��݊��#��#��Л4�+-ݎ:R�����������y�uP��-4Q�_��XN�z�\5,�1r%�I�&���������f�Ca���]4
<���ԥ2$eCg��$�nu$��lM��"3�!��v����x�q� {n;��B�3f?]�s�+�V���L!� �K2
���QUvJ�>�2 �Ӎ9����҅�� ��<gi�'Q���P7y��6$��<y�[X����(�.���_�(x���:d�d���&C�i��@��[D��4��j����XIG�٘���&�Uq�fv%���]�(�}���7?�K2i��.&�!l4��˽�6�_�܀���f�[|�v�o��N�m8C����iLR�E����ʂp԰���٬�T��[R�=��)� J�Q��/j]$cK��Z��Z�7��`T�"ѻ5�d��WN"�I�&��A���F���ϫ��b�F��BYޟ|��G9`V��}V��|��Q�'N�Y�%�t��Wŋ����	T9�������of���h�!��RE�@}��{yS MKDwet�=ȡ�i��%%}�n75��Hֿ