XlxV64EB    17f7     9b0��b�O�� ��z������6�-L����P�+(�;I�-�ͼs��|�E�XpH:�#��v�I���R�§J ;DED�H1��YB&Kȱ]���%�l+�x ��)@Lw��P����~j���G�S�N� q�|�㏽�·���j�椦g�����Q�	DŎ|�������ލ=�A)a��=v��s��3,�m#����j�LEd�U�yH>eRz�u��N~yjUϲ4�jV>Y��f˝���PW�^�)�V�����j���Jǽ��<���*�t��pB�ݢ⚨��h���L}�B_��x�h`]<d�_������`�u��C��	��o�?�a�DC��@�w�����,�Dŋ����˭�5V��V��I�C����&Sq r�>�r��!��t�T:ŋ�����6��5�F�7�	m��%�QS\�a��n�ܻ�Usp�Bݯ�h���O���R��AE��Y~��X���y2�͆�����)I`�`�-����GJ+4z]��|׶�H�����-9��1��h���	�����/���ػiab.A��wTc2�����Ž����=țn�Ts?[xɛp�}�uՎ�0L�h̦#Q+~������2R�RI*=M0�hY��)�<R}[Z���Xe�X���	l+2���.���fnu�C��1��({r)�r�j�4 ,\kP�J��83�D�lf��~Vgjp)l�qz�ݠ(������J�ވ3+r��u�S-�a�A��)]��A,!��D�o!�*�(�G�j��&�$�ZCXC�~#Q\��UEO���Pt۳� �mfz�xp�=~5�l���l>�}5�1ץ�T�L��Ĭ�����,�(�_���c�������D~�G�9�Y�m�A����̩i�����L�Y�Ǧ���<�L0�x졙 D�����\�ͼ/i�*�(:�A_�����9Z���T��`O apF��Y������t8�f1��,:m��ز���%�l�k����I���^�a��l����A�L}�sZ�K�Ӌ����\�	-���[����1����#I�C۶����I�j�O�%��c'Vi������A�%���� �Z̛s1��jlF�yp���ռ�rL�yz�ݥU9�ё�1�����d�����x�=NP�u�WC����Y���9?"���GUϞ�}S�������G`@yI���tZ �̡���l��"��譑C�è7�C��4�*ȭ,�G]�$&��+%���'�C�ڙ��r��F�K]�q)�P��(�+���,�/�.�u�\�>�@�+�ơO����.���)Ы�lr�#�����;��q ��s�3w�	@��Ń9������y�?��c�:���˻���Ä�.ވ�%X��&E�'�\@Dw���C��E�D�n�>ʈ$ZW��F�S�H$�����6Fڷ�E}���,I��S�N�^�|)�N���� �-��p� -W�|�/���HV�(M��L���m��#Q��ʮo�E��������̖�����%�3���}΍�yrDI��}1B��	���6>`:���|�Q��lᰮ�
9ɭ^?��.1�G���z׊S���%e��������W<z����I/�;��|�g���p~���������,���Sa
����dT����
����@Ø�^%|�Yk��x��D��El^y-+^7�&>;/<v���\�����M������%ե�KK|�	�\/�qZ����B�K� �E�z��ɝV~�ey��x��1@�Ƭ��־����d���]b�P�֞�$|�u^�OS�.�^�H�=�jŞ��+#{�P=��w	_	 r� {�B��Тʖ���b��OHy�Tyݱw�P,�c�PĞj����	CI��e���1}vR��yr	L��e,m���I�
o8��k�����	:;��q�8����r.I�cᰞ;���7���AԠTc�x�?���9�7K�z�H��Ϝ`���jv�ϯ��&�H�u���*�1ygV�r�ėV[��ѯ��}���CXH��S���m�K8��M�G�r6zn.?^ş��L��߂i�-�)<gi��f���y2����M����*~�%���c�efH�&����S�ه5�����v9�/�(T�r$%H�ZL��[
̢�8p��1�{�ұ�1���z�בh_���*��D��z���"�fw�W��PK[̷�n43�@y���*�΃��$ ��VՉ"�YOc�@;������tz��R�~Θ���	��Ɲ�]%ݧ��[ L�
��!Na[a�k��D� �����4]�J2Ɔ`VB�V)9%ɝ��-�����GJɈ8b�#L��9�{��A�uιVF�U9���vA
��,B.�tr�N�#	&��So���x�?N��te?�����q.)�\!�{�t