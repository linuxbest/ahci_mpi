XlxV64EB    618d    14b0�\ׄP�8���'�%�+� ��G���&�� V)X��b>a-�z�`�azDQ��p�&���z���}�3�j���D�}L�E8'��"���EerFM�������!i����
L�	�t�����������)�\�V�w�o�Ι�I�p�Qa�h�ݫ�����ڈ�C.�VF�c����z,f(��HYG�!i6'Q5����C�e�2~��3e���Ј�0�"��y[�׾Xd���D���&���"��Ngȅi���h/�9�q�'�';������mk�ː���q�����?�<��NkȀk�*t��i��RA�Б���pi��b�"�P�@*�8�U'�G�z��jɍF�+-�~+�y����_r�iz���R
�5V̨��ϲ>o��W��C,�s��a���j�oV9��&����{��e&y�
j4��O)1k�^irn���e�{�[��-����l	�f?����I"��\����i�1��6j��ϝ+�#P�,��D��8Y�36�ΕaN�K\��	�]���6��vf�[�b���NYsԧ�$ #��~!�%)"��W\%r�XpY�f��|�d��������������%̊��;*�פ�?(G����)7��G4�>46J�Q���p�1Z}�t*m;����P���'ۻ1��F�}������	A߸�@ ��,:���z�D��LW*m�t����AlJe� 9Z���c�U):���#��-���t��*�s�CaҩA5���5����G�P�Vp�U�N�&��� �|t.��'���؍be�}��;]�z�4�SԳܷ����T�)�d�: [.��RýmRoAxW��e���6��8TͰ;�z�dg~5YN'�M���.`���U�����s��6�m<|�o>�M먯�݆���q?u�<�����z���0C����4��$`k5W1���A����Ž=3+?s
�@ԉB�<���~���!1��. +;���[|�3��T�����vЬ��|ɢ�
��/e[t7|'�i[)���a�m��hZ����̥ڮ�FB����}W� (�npR���P�:@�����g��jε�t^z[�L���xC�◤�m��jI����//b =-�`�$Hq�N�X>��.	*0�� ����-4ρ�İ'tz�Z'����W��p��j���;5.�����L��ǘ|��9K�Q���0fy���T��IZ��r-�k�A���K3������8Xt|�5bv垴��	�&z���I�]��5�ˆФ������u���%ݶ�sp�Y^�D��ù�Ս�M�4����3�i� �8
�E����Ҽ�Z� b���Dx��#��Os|!�z	k�h���ԗ�_��󭎲��z��ng���d���%j�K�kF���~��Z(7.#���b���H$�? K?F'���[Fg���g��X*��������������`<���C�7%8y�����vs��6����s�s���Dy���(~I�G��Y�s��he���c%�:��	1$sM'u�H�����$��/�)ڐ]�"l�G����NV�����zs_�����w�ü�Eb���W1ΈR�-!�)���vD��7��=�^]r-����*<P���j�3%������槳�\�vY�T���d�4�<*IV��i��9�EF�6��`ޜ������h�lA�	4O�#Z�3m�\�Y��_��z�㼡)>�������$Z��:��z���CZ(d�`ͦr��TBm�s`_�k8h�@��m��D*ӿ��A�4���9q~B�ǈx�q��R��S��n��Ĳob3
Pűub����G�p���H7�l��*����|�	X������C�.y��ϾP�ˊ>���wG�_�
�Ƚ�t���n`V��0�'һ��W��ȫN�����|�h�~����{�F��t��A7�T7�9�A���;ԭ�^ɮ��gI�	e�Z2A�,ǘ�S�%ۊ�����몟"o-��	�tOy�o�K���0S^D�����v���+W��w,��<�u��
�1G�)E&8zBa7�G� 1W�g���/sTg-h9�h�mB�%W�ҳ+'z )�B�n�M�V��<u=f@�y"m��8������e��T�Dc6J�3T�^�d\��3%N�YRP'�џ~���+���y�F�+K�m�=,�Ay������V`�l7�M���H���>�]��*��:D��׭�6�ڣ�����3��Y��ue���+:u�X�D��]��&Ћrø�˝�bv{^� ��R��IDRV�;���"��c��f���p�:y�|��f�&�\Ԥ�tTp�1��g|rPȜe��fFz�Z�A���͊�lg��s�0�}Mh�`a9ˤ�V�\���%�H�#�o�Bվ!�~�~7(��.�r����b�����z��Z�lE[�D6��!8Vm�L�����G�L���Y�2c%������3�Z�SV/���L��J�D��A㷸�֞#&�L[�0��s
��NI.	y����s?�|s�\a�v�PN�f���������{�SI�K�w,�v���bd��u/.�5aM�%�NƥL?�<�0M��7+�'����{o-�<J�G��Ed�
���o������B;�X�:/?D&����_O�{��� �T��\c�kH����z`_�\�wfP�{������q�02*��sHҹ&S},̷��3"�e��@$�nB�L����p�N_�78��a\�)Ӡz�����Sd�o�#��a)I9ؘ�����!W�FM~�s6w�&���=�v��\�5��L�^⍭�3���r�
���N<�>���[�;{��#˷�B�k�!h�_�]TMW��(����2j��rp[�asY��Y��VZ�垆����g�p����z?��q)Iΰ��H��Q]݁{��s��W�	���֚�C��!?�"��_xW=<�\�K�f��K�
��؞�����p��E�شɚA$nd�(�E��*�;_��l��|�p����z��Zy�M��&�E��:��c��%ZD�S}1B׺��ߦm�O�ozU�F�s{����>�ձ�fA�D@<��n"'��9v�)���ը����o�E���b���~�����YW�[�E��|*exৢ^m�h#��:Q.
�^F_����Hm�:EG9�^�.���G?4$Fm�h��1J3NW��Vd�s5��PDH(�).�eȮ`� �������´O��}�F:&��C7B�3K�b����!ح�^�?B��\`��g1^�o�iG�Ԅ7ataH�Hkum����=��1��!�^�,z[�Q�A�NH����v���C�Vl�y=�C�Ob��ľ��~g�F��}�.YbKO&C�����p@��4!^V1�B%�0ِ1(HE�p%�t
��e,w�]qK�ek��tB��.n�E�*��p��N��d�%ؿr���OQ��B�'bc������rĤ�=ō��-8I)cF�`2,�{�!b=�J��+�U���Ae�6��{���Q�5^F���9�!m2�U{~��B�Ϯ�m�;a�p]������d]&ak���|`l��^i������zr�7 ��a3�`ثk�t�H >�}�\t�^䮽�%N[h#s�2Z�Z5[b��Җw5���d�mQu����{����1:275�xWw��q�D�9����`|:qoH�g���u,�d��q*eܨ�*]}�����Q]�s?]<��AoN�Ir�I_jе�b�ȳ�u�<w�����MdbǺu���c��TŇ���"��h�L���?�|'�Jy�O��Ԥwi�J���*f�M��V��~�PВ��*��kR��<XY�c�����Wn��{�oiMR�"�N���zSP���gV�AN{��>8�}�p�Z)�e��׼.s�!AIpR���xg`���?�O�����%�L��	��n�a�O���6-��-��=N�ox��	�63	�,�zDUUM~�J-Sb�#���9�/��Po�
��I�^R5��@�'u儆q)�r���H��!ܗONMy��o��F�L�����3 bH��Պe�ĳ������	c��A�Y�z~�.�B)h�3�vw���N���c]W���da�ُ�ܞ�g�ݮ�������חP�6;λK����,����P���x*1�I1Nf��d3����i�믈}b�ϖp]�S��-#�tC�p�v� �`�G����f����V�{��/h���(	�f ���b�x i�g�i�4q�
�dg���cXV[)(�@D����3f;3e���T,Foi��u0S^!۟\��d�
�T\�ب��<�[�:@��G �Ug'mbd�!;��n���s��ĺ�j��D�KgU�B��#��{�?G	��@���`���6��Q�i��>�)�'���9���'hy���C+��>�K��Rٹ������2SLEN����[u�Jc�J/~օ=�u�6��*�"�.2	�0��k�n"�!�`*Q�k.�r;H��gH%�Q��z�5��S*_�����GOS�p
��b�e:,�̙��ڸ��a�7YZ����J^y�;�{���H��B's|�I���U\�墁<�J]���>p���1�g�r�B9���쭀
Du�'�ŗ�����
�noR���s���0Ĉ�!�jH�E[E��c��`$�B=�Ꮕ~����(��xO�H�I����eeru�CtA$QA��|�!�kJl�����g$e���ۜٔ�K��Q��W"C�����]a��	�/���O�5�\�1E{=�������ǆ�-,\�7Zq�1���Ͳu��.��PJ�PZ�-�?ep�����f#y��1�ݯ�Գ/>b����P@If1�"�ETk���/þ���!\�ݚ ��R����O<m9 s�aAٴ|)7�s҂۴����U���z��f9�=��F��x���z�U�1�|Pb2%��C��f�*5'���	��n)�x�x\��5�P��+�����h�2�D}�фG٢��)�)"���SK�5�2!ӛ���2���:	��cS����V�Lv�g��dM;'��l��/�y���Oiz���q��.��"�Ҟ��"��Z�	����3E��d|S(��3�.�Q?��@�A���	��vJ6_#���f�e�c�I:ۺN�