XlxV64EB    410b     dd0G�؃A5�;I�k�a2.8h~^��7�E�t�'�q!+x�'�VM��Wf[�ĪN��^Ӳ����
ԝ��B����f.���yq�{6�Cr�����=���uME��2�dhS��bx-yB�:�?�yuuAE�)�@�[�)�gԎ+��`�̺�[�J�S�mmg-�`�8p��ʩ�<��ᮮo��a��D��C��2'Ɨ�k��B>T8�s�d���Z�=~g�t�篱ۄ`�^�v�,�D?�(�͍E��In�e<�U�^Ou	�gɛ���`Ҡ{K�*�����e���܈�f^W�Qa�X员s��p��I�z�@�G�I'���Q�H
!i��1��F9=ʀ
>ɳ����g�
�U��*��c6�h��|��Y
�9������OPR
=�K�3��c%��aCUJHs�*�����_�0u-�qjE��Y���Z��(Z�Rua�ÐE	�p����+Z�� z�����[0��2��a��+�TiR@y-�]���Ġ�U��
��szĦC]2蓲�R�ZfV�G�i�<�� �5�� E�v��D��hs�O��u��B_GNzz��&��� q�d2�Bv�O)F�E7�8�t�%��0I�@�Z��X�� a����5ES����F�h��;��%����p�=t)2�] �L�b�'����Bi���In[8�0�DuҀ7բ}i-�l�K���P�5�*MW���	��bSY���௽���s]��P%��^]ؐo�Di��=#�A������Ѥ�Ar�t��4�?q3��2!?B"Wu`�RD�%��{U�N� �z�xq��[1U���l�7��5���\r�n+��?9��l�֧=��N[��;�����<�Ld���t]�L�&��ps�wG����x5"�$��rgvEr笒��j�F��Ň��8�A�!��ʬ#�Y3�a6=�n�±Cg�u��a��N3�,W͂S�I�c�fu=�W�����Z2辙@�����l��R�uj��<j7�	}�8ؽ9�*f���Ge��X%b���Ѻ�O/���|gw�D��
)n�'�RAD�QV�Q�4f��y���~9�V}���X�_/�\�Y�%�E�x���h���*�����tɇ�-���B׆$�_����seQ��+�X?�L&J�{ݧ��E�ˊYΐ3z�j��C4���4��n�;0^�.h�E��9��w�t����V~�a#=�䙏�C�S�%q��EP��P��0t�A /�/zg�{u��9!�8yQ���iI;#�s���D?o')ogT��������ŏ���6��յǶ�"�j;?�>ÓPej�O�tzv�/@eJ���FmE�ˢ��c�o�@h�KP��9|wE_����l�y�Q`X���jB������P`�U�O�_�U�/�$w^�����"f��R��.e���(3<�8z�LD;M�^��m����`PE�,��F�7p�Z&*�'G�ڶ*)���D'�N��9��º����g�~�뒉oS<��BC�B_�{n�޴��9�t������̼�$�imSh�����@\�f���7H�Y(Top'��_]%�Tk9:*|Wf�)�t�-:f���:�
ZB��
=�����P��#��'��.cO
�WI5C���;լ�7O,H�{�"qM��$����V���q�)p�2�s�0Y��AЂ_u�����%�3Ny;t��%��w�؄���Dz4RTP���J�^h�Wx� s�Ώ�j�`+S��h �v���~�A,=�!����)�^:��o�����>����8/��A�c̨�U���-&���t���$��e@1��:��y�oe{�;0��@I@�����ΰ>8���hS!�ƻ�R�TL�F�o���{C.P����m������5"Uĳ0�֥B�6�J���@��\S��MH�1i.�S�d��+���0�TԱ �i'�䷀�ဆW���*�q3'Spɔ��dgAφ:�D��dfD�{9�Л�Q�7�M	sh'T���Hs�nzR�c�Q<l��}�!^�#"_h�F�Ő� �UZ��6,��pru*�K(`�����ةa��9%MAx�����a��=�C2i�0�g�vu��i?@��j��6{
H���V�B7�WRB!�r���#?�����+x⬈����&�m(�2����l1�j�F�y�cMN�0}oȆ�}l2 N�s;^��:4����.:�U���!Of���а+�H'��J�����C	�(���[��ܞ��5I;'�[Ta�'[�Q+A��Z��ZN���냵����H �o�j
�AS�x����� ��BG��@�)Ll�����u�Ene��aaW��A�5f�_�B��
�-Y��Idc��kUQ�
��Dmq ���� �c�ī�s�c�F� ���]�_��*Q,l"� �b�pe]����l�X��DI"�	�O�/��P�@
��\k����X��v��o$9������zγ����:̒���✱U*7� �'�����_@Qb����Ia<�P�l����W��i7����W1I��-�8�h%h���m�,� ��4B�K��̶�,�"�}Ë@O�������~��Q2�E
��ءz�QU�����V�T#�W�eCPe�B�=��ךm7�m�|���|AyxZ�ȵ�aa������t-T��pn's�6�Ģ��0m0��)�!KD\cI[)�<�����uHjs���_k��yY��[<�����&�@��O�OY��l��r���jQ ���ϸ{���gc���*��u����"�R�Oa���9=�,�Ϗ �.��,Ft�@�}� �<�҇���_�&�f_��)W,�+��2h jڛ`%�3!3�WL2��?��Ț�䝡�k���a�:9��J~Ap3p�f���X�S������
�tGbߚ�$�4gBK��jq2Ov����j/w�t�V��W��-�z��7��]M5�S��+�p��뇲��O1����:�j� �Γ}~���¨��,��
�R8/~���l� ��K,�1.(r#��AT�^�!@XJl^O��m��Y��~�!�~�*�MK`�,�9'�i�77(c�T�
\� �U�W�׆�b �/��>Jˬ�.��./�(�c�{��
���g���+��q/9������:�`+�;E���?)_�?Ŋ�z���/��͵6N�޸M�M��z.���-3�B1L�kÅE�P=���~��H�?\��瓵+��t���˺�����M��<��!��3����{X����zS������CvI�?V����E�9įy���K`C+�ТWĭ;�I�SY5Oq�$\�p��3��0H��\x��� ��D RF���U6���V� Lx��T�%˪��9�@j3��H�D��'�VEEC!��cR��hr��[�ܪXj��3\�uJ� �c�&L]Ҥ8��ڧg�����XC(�U�cp�nU-&:��ƕ��p���F����