XlxV64EB    211d     a70�+�qɗ�5��}���?����-�ZZRÇR��+��L�����e��q�r$�k�����7"lx�,�ud��k�!l����������4��D�!rl���!�,3s]�Jυ9�
�v��E�Z��h&�ػ Ƈ{apQ?�3ϙ�J��'D���QG�d�}sdS���I��<�ͱ5�#}�U8lZj���]�?_����b�W�qjeUa.C�An��N	��C�;��E��_=���1Oz���A����#Y�wh	51�X���iU'U۫h�d���`�qI�zT�l9�ۉ:���\�Z �:�Z�:���()���m<�.f�B�R�涟�/�H��['y�H��;CO�8'� BZ�*NRj��O��¸�*�̉o&']���X�c�hu�R�ѕf�ӱ�������?������2��8��fG)�e��3Dw�?��c��5�?]i�΄���)ظ��
IN���;3��v��O��ˏ��J@y������vkq);{z+��㚱Yr�ԂHu'��xN��QԨ�"�#-�*��u8Έ��'e���&�"Q��3�a�Q��+����^rhjls{a⮐̹����%eT��sLc�yz}%��|��W����|�l҂�3�uv���37���x��t��]�����Pe:K���8�P��݌���ݍ ��}�kw,chr�Ct����<���[V��t��P%0F�h�(��j��$�u��$Q��3%vmb��*4y�H�$��g�U���� bρx��K�>�#�D����PTCz�+g�2G�����xN�'c�|{�r�$|6IԬXo�:Ʊ��H�T컡��4�|�����SuBwLAV�JX���X�^I�R�Q���:�ػ�^>��xN�7g�f�/ԇ���8C�e/d�t4%z	��R*�y��̉+�m�11!�"j����[�*!����qt�K�:��W���YǕ{C/�&+�g3_S%��s���d��q�1eA��k�E�X
j��}�G���P2�GT���>���C�7QyL)ڇ���]diYp4#ҞEЦ��Ǹ�o��=�>� �T�\���)y�3�	�^}'|2|0Pq��f�p=mYE��E�ٞ"�ߔn�S�J��.e��l��K���X]L�#ϴr@��@tF���"q����DUb��l]����%�9�T�sk�t�mK2�Tۃ�M���>\Q�EX������ʏ+�t�x�+�0�����n��"}�A�^�C��,=�s�o܋��1Wׇ�����[�E���(�쵥H,�#r���Y�.��t0�w����oA����C���AV?���\����E�ũ��LM�[m�,��s|��pZ�� '�Fb�WuV�3W�	�ܒ]i��Y	�X;"Jk QI�-�R^��nfꊋo����o ���sǊ�[Ya�_6U���^�=e����ã�����SזzȰ�^f��$0`�;�6��cbB��ίN�̔��i�6O�Z�_О����v)�fYO��V���b�U%1X2���k��bW��@�O�^��|��n>������
Jl�ta�����x�.����w̉,��?s��[�4d.!���K� ����D@J���:w�@�y;�1�����0����)�B]��z0_����1�I�y��E?�r������ؙ��؍3#�2��u%?��T)�yWIw}��Ļ�#A:�yr]�_�:���t���(pT���eeVFw5�;|DXq��O�r����5�ѶeB��]
��#�_m��:��W'5}x��^je��E3s�f)M���0��Z":q�d~����5�����\vdT�BHq#�����`�pZ�Q����O�E��LD�#�v�9�����`]9����x&������Ӛ�F\�Q�@�G�a�?�� ���S�|�������|������ݯ���x�|�`��sIࣸD�
�)У^k3��&����EO���j.]���r��mhoa1>��Dg��������]-�-�U�0�p??n�9����T�q9�c��{~���za�R��"YMė^dg?^��:���!)�ȍ3l��^��DTԆU�ĕӣ:}��FL��5��wT_h�o���L@ϑC�,#}-w 8~����M^��W����̙g�蹡��2+�vq���V��0�U�L-ڿ�ҟv�-:�0! t�'�����d�;��"���$�a�N�z��#��GSf����D�U�xRd^��Xn2Q���bgo#3���[�Щ[I�R5R��^k�YHi����E��ʪ�2�İ"5>�_*&zh��%u��� ��2��ݚ�Y�+����M�����qQ��sh}z��D�rc�2�o��]e�X�M3]M0O��D��9ѐ?��:��<y&/3� ����׌�ڸ���'V�G�8���e6ͺ����	����'�۲<�>���ݛ�f\TC'>h�u���}�o��NH%|#~�8QM���#�����k"��	�No��A�E���a�x���jW�웲c��v�+O���u끆��e��U��6��X��՞�"�(>Pm<K��0E����I")���f�#a+�ywv�D���Y��L"�*�QUw�j�%���k�7�|�x�$.1�֋~���`��*q��V��JUb��/