XlxV64EB    1b93     9e0��a'�"_�j	�m���uP{ \e�Z[x����5���"`(���t��V�a1{_��֍���&}{��`���ZX�io]R�Qe�$�hI9{��h*�!I��w�F|-��ϼ q��$M�'�[ً����^i~�.����\'�9��ҝ ���.�e������(��7�ѮJR��t\X5:dxߓv��Ή=ﵬsh�Y,]kV�U�`���~��xG+�t��L��+���1�ʠ�:+�ԡ�GS�[�5���<R��.	G-[�@�M{{.x��
�О{y�m����ET��
�c*wl�-�	~o���k��܎~��|u�UU�
ܸ��gn��}�
��$�e�����=��<�n��-x2]��,?��A��TgW�G��WY�����8H�/����Qp���|�'��1����ǀ�Ђl��n���i�2����IO��&��_Sp$�i\J�z�i��Z��y��r`�)rb#_ӫf7�:	��>�}���g@;�h���zع��?�6\d> �m1�t�oh�����ۗ�Y�E�|>��U�Z�2�`������D�~��I��aU���ޡ����}H��+�&�����7�jı�X=e����G��#1R��e4ﱮ�]Ś_�=-ÆM9�IQ`�Cy����ư�q�dF�p����D�0&w��'��tym����(��[	�Cr\�cx�>��[�+�NN��ΔJ*�4���U�'��D�ݗ�wU�f�^'����Bc\��ݦ�(pqI��#�����8��z����f��n���W9��E���MH�g>AL4�����$CSn�2���!K���+�p��"G�������\]xb�>��!��b=���(g��3�WD]�$؊��}������7��T�ޗ��m��j�@�=q\�e��H��t���	&fI�k��_;QՁ��#����&��/�q�6�9������E+�n������`��UAz��\q�R�ˠ�#����t���n��>��q����{�����Z��'# o�3 ��v5�ŉwS c���>��͋����b�I�U/����coB���Zf���f�|;
��5��:͚<!Ut�6�YZ��Ls���z������[D�m��Y��h�f��a��?`�a��cJP|�&} �J�_�>P�{�?�l§`K�� �A����Ț�e��AQu&L��/7؛^�o���
y�Ⱥ�Tzz���~	RJߤ	�q5��i��BFu��>��>r���g������48��1�i��r�}݇Dz�kcK�m�_����@�Y��+`͌�慱 a�ڪ�3j>��!Y.�?:�*<u��s(Bm�#L����.���?m1�c�&�䁐�_���߭)R�3����B&�E3����I��K��\H��P���#y�h���V���l��u��Ixi'��r0�+K<hi���$������3t�č���$�,!�l����I��n�T������ț��.W�ةO�`������7g�aüN߹L����R1�\6�nXp������72_,#Pf]n��v2��ndV���˧��m���M�#=��������A,M�GY�g
$Xք��%����� X��b{�7��#�9]1X+���+��/ŘR�vq)`�����=c�"���

E������c�#<L�{���M2ǧ vDw�=t�/ZWg&��{VkDJ�1��~�$F����nd!�U�Bc����+�1f�a,�EE�����G���=a2aHFy�n�4>��v�$����/�W�h���Zѻ�K����m����_*����u�n.Z,�Ybs�>\�5:m-��}i�5�H�h�N3�i���u�G|".��|F�,yzR�%5��͸�j'�����+��_,�_c��Ee�e�`�A C����>?����h\���g�q�+bJ�'G&�����͍�x��v��>�H�~��P[<�f���q��J�w�[�r��,tB�@��$��Ә�9&�4XM���)J�Ͼ����cQ<_5$� ���&Il3�+lqlj���(�NC���r�WfN�Nx��z��D[X�߰�o�hWc}�구�g�3~l�J��r@�.0~��"�t~����E)�	 �;*�L!|6�v��������^���M=*����ǘ���k�3i[����h�G`}����@�t����d3f�ǌԎ�V�E�`��Z��U�M����Q��XG-�4iH��{�� &]b������;�|����蟖G\�'�k����k�.@�w�KZ����{�>�JƲ��w�i����{�
����4m����5��q��
�@Ad�D�N�h�%;&a��J =��?%��J<�`i�����=<����.M*��'��/�P���6�Zw"���&c�-/��*���_���:
�4 �t�����>�0
�3b0