XlxV64EB    9710    1dc0�z'0hSu#�>���t��l�v.����Y=�n����煉��q:`�� xc���-��H=!t��҈{0#9T���o L�Q���L`10�8�ߋ0�(. 6������\� ۧ�z��Н>r�E(#T�t����%�>��!a]�ZM�|��-���s9����7�sȃ��nU�12�f1��c(�ɂxa޿���qHׯ3�w:؟�Fo�J�F]����Uj�9K�o�|PX\D�g��/�N��c�?ja��;kDxŌ\��fK����k\5�+f��	2�d�A{=Ip���R�����hm�C��7�!�(+n���4��v@aw	5d��V1�fjŞ���T� �8�%_Ӕ0�eM��$ �ф���CT7�Op�()���E)�t���W?�Ο��Y����j�#���b�B@�v��h�wڍ���CyA���Z���ޗ��AÝB�6�k���H/��W;%������,wL�=����P��rhNL�g��U*Z?�Ei�rce�r/�+_Ä�G��/-�ٽ��d����PL�/Qҝ�[����Ⱦh�+"���-Ӄܜ0�6u�8�A�њq�3P ��Ԧ�$�`8�7�b��EV:�]t�D]��y��]�H���5@��x����{��JC8P;9 �����Jw67?8��8��_�~軯�k/.V�2r sp8�5��ѳ0AwU�Vc�؜���/ �+t>¸A���E���V���_7y������"�&;��[d#i��T�/PJ^��c�&E&�_;-�i�_���S�M+S��D��J��0hR�'����5l���������c�Ķ�����8ax9�´g��m1ym�Zs<�J������u}�߷�XNёuL&Um�
V�����K䝍�%��k�2�Ǎ��;�J揬��#�M�q�������V��᫐gCc�^����o�~0�~4(In�86c��n�W��"~uޤ����p#5#ImT�z:�Zaސ'��!�w��Y��a������]��)���{r��AGz�/�'�z{�}jaK�}ec���M'ѿ,�.��v�X��j�yp:�#��BEA�g�~yWHb*-��V�!����ѿ���/?�cI ����Ŏ��dɮ�z�G���g,-v�>�g�<����`u��{�]����W��� 8��f�V Զt���W�����$G�ԕ����r!��5�EHHZ�'�ע�h��k��P��Vo�.T�.��LT\��������U�o��K7�z<xg��1*S[H㨾s�6g0�Ծs�G(��,��-	l0� ��"�"ؑ�Ȕ�8
�p9�<e�:��^n7��!1\7$A��j��f�b�ڣ�Q�HY�w�<`;U�9�2�'���W�d�@��E[Jw�q���SK5�q�:�uU������.��;���(}���{A,B��icV�pbu^:��t� �L����E�����P�� ���,@��A,���`�	�xRYo.�J0�\�T�_�7�}Djw�ih�H�]�/>�E���/U�||��Of��f��xl�/��j|�}��ĸ�NlS���}�nh�g����k�iOOE^�+SQ6^S���{/���Z�K?�T�\�<쀋�(忝�k}�Z����z
6t*B@���J�+�98�~W�Ҭ�*�7N�A�̜�3pkH��G[<�s�Ҡ�D�����A�[>&���C9dE4\@iTy�$��<;�9�����G(�&����� rO5�/��QZ}<�7�Y��?΋�r0�t �W�`��w�F�cB4e��1��I�n'I�
7��qE?h���U�`1����0~�*���-Eլ߂��,oKBg~~�Mվ��`>�w�j���Vnz����%�)������;�Q�iK�[�Z;�����a����.�9�g�P���7��-m������@�IFgn�������W��4C#Ю�R�Ok�졔	���w�;HS
�7���h+��@I�:�ڋ�Qf�p��бH���.V��R웙x��G��MB��RÌ�E-O��s��oUj�8p8f���V�G3�����B�<�AI�.y��h�9z�r�}���ӪQ���=�s�ɪ��'�i�s����� �:b�Jt������Kg�ďE#1�.>��%�{�)*2&{�A����1l���Mvu�]���b��}5{�9�c�&=]��>I�|X���_��!�ؗJ�Z8z`L���Bf�cRgשOPq�YU)��ǫY����#D @tW:ҥ�_��|�~�џ��1��$��y�� H?���1���>��Qz�$�/"��)l����F�F�ن��i��m��^p{]�.=���;o���)��J�s�p�l7������
����(�"e����=��V���V�WT[~\��w-�8���w��,��O7wi�I�z��~�Db�φfʴ&ME�_x'�;9���G$�[IE��^�9V�p���߃<�r��A�j`��S���ƙ7-��a�w�a�]!#�T@Wa�(��G1v�ĥ�4��_]D��f�!����(k�O��� ���!*ށ��Q�����C��EV��wv	Ս�f�"�}N�ѩ�L���Tx�>���@�C�Vc~'����
d9�6�\]�U��ER?^���]���8U���Z��q����fa�UdO0���IDd����Zj��r��8ց-�S����'��f����b�N��:�ᮥ��i�!��u8����\�XK+�+�CL�������.��ENB�����>�v;lb���Zx;7G��>\��|T�[~��M�)���^����~��ɺ����[a!��UI��� Nm��Tmh��wh+Ap[��,���nt�!<t�����hJ[����?��>790(�m*��`Z�?9I��L1��k^���^'���o('�{N���@�=n��;���X6z�:Y��:OڕK�^������\[rN�'�6?sr�[�7��L�4e�}�������8SwW��F�Z������e��r����K�M�/��[͸I_n���a
���g4�%>j���hl�����]��Ĥq�%H\Rf�F����*Sh��QLaܯ�w�ؐ������)1?[@Oٿ������^iړE��BS)���e�!�|ޖ��HD�5Qw0@�D!ٽ��[d�L[��G.�kƋ�"%Bp����X@q�D��Yxn��ˣ�N9�^2�6�%ꢢv��z�c�	{h���|�g{/-��L������4��H����0y3�����h�U������A���>�DPl��=�N��a^�"�=����^d*��ıǰ���5.�Y�����k����*�9�s��a����J����l]jZtK��ӷ�zJ��4�����R[2�mR4�I|�o[�Il�\��u�	�����|7�s����i��a���.!D�L��K{�k��F❜��?�S����ΰ�d��ҋ ]v����J���|s���k/O6��l����n��g����@)x��Q�暇�0��rpQuܥ�x�-2p|$�i��~)j�n8k�)߻���2/��I��J�-f�9�T�L�t"snc����E����vnA��Sx������V�0L�M�����؍�v۫��
��~�J.�h#4Pv���9J�X<j��/(�\����X���/�F,,�aخ������o�\���ub����ΰ���9|I�̎������<u���J�:<��z��l�ywP����dy�{,d��r�2	�
��;~�-��U�4�!�`��Q�(�yXV��'���M�	��K�����"�̯=ˇ�� _a��S�\�j���5��3�=�}�(����'��~9�ct�Ԣ& kxW�����QB��VY���f�a����6A�}Ya�r�V�/Z S���c~U1�G��8 k��5�w���f�i��x`�-i ���r���'*�Ό(N
���������㇂@&�zltKxz�g`@@!�f���治��m	6My�^E�c��N����#\�?!���P[�����+��.���O��\x��R�N��D�-:�}3��A��O�s86�Ub�:�����w˖�p�zA��$��6���]6�1���
g��Q�xk)���Au.>�ePYhW���:�Bc� �[�g��s�|~epW���%���1�ň\����ZZ��V7zf� ��W<3�i�8A��=���km�
o��Q�r��<�~��d���:*�����˼UJ���/T�m�Ł
�)A����)y���0qG�w0�������t����!s���_�\��4�\���Gb� $ف������`L�nntfO.��<E?�����z�������O��˚*�%X�����aX�K�X��o����b��I�Qu�Ѱ�DDjL�,���X�8�iN�ً����˓21�,���Q�&�ϖ�s�?}��'�	��F����͆�0)A9�����Ys�m�����Vmd�WR�^!��$�Z��D��U�;{�;�qS�GR�{�Ó<?��$�/��42
�|u�D�QB12�� o+D<�v��uW	�*��in��t�X24�e�9͞/ ��[ݏ�+2��ú�A�P���/.	�nW� ��8/q�A�:E��Qv낮0�A�MѠ�/�����¦�����
{�Թ�����u1�s(��|�����s�2g"f@�|�cH�n�^p�<�?�"����v�TX����۟/�@L^����BJ��\|^�<߻\����۷XV�>������mu�įT�7#���6+�+7ѭ�#t��=��XF4�n����2�����K�<`�����J���<ـ�4��A����6ߌS��lr����^� Z�%�-aσ���pd �9,c�ő��ŉ�G�C�"{�����z&��?��y��}�5R����tݝ&XNCG��F��Dz��jh���H>|�$�m�HS� �Ql��I�>h`��� �@�̾���N�'@RO%u����6��2;���+�>-B�RR&n�3/��X�+`��X���XJi��[�~5�sK�X���;bHQ�'yLE@��hH���Yz0�f��&J::y��D!v2��z:�������!\$��l����&���,OK���_6�O+�{Q�b��{�O|%�p���+:�w��֎x�Z���V��L��iP�Pe�dx"V*��]��X��/ؽxA{���O]e�S
�O�?���E����:?��~�Oɗ��D���",0,�&	6X�I  ��j$�w�����#x[w[ӽ�j�a~��lAqb\��#���?#0ZvZ�j�0q����EE�K���`����W�swH��%� �̹�p��sc�=��&\嶧��3�c�Lk
�QW	Q���^���2m��q���ܩ�NPtia6v/N���&�5P��(�����e��,fXx�C�wEa.���&Hk쫢��v}��,n��."����UZ"�ҿP��E,���h����S$+*��>�O ����2�0���!�u:����$�'4�����m/���"��4#끍���h>�Yw6�M7�[�5���A�ǲ�d�Ƙ����>��`,�&��=�P3�o�_>�ٽ`�b���m˯����2�v�/��2�8Rj���l^f`���ZI�a���܎��HO��⎫�.5�2q3|||Z���RI�q������)S�mҥ�x�P�%��M��uo]� �g�&xB��t+{2ƌv��g)T�Wt4Y�V�Z�e���n|�Oh�+���'@��MՎF?x4H)A��C���
��G�?�-���	�����?:m�~�u�MgeQ�t�_�`P��WR�%��e�y�$�e�w<����d����j���|��Pm%恼L(IRk��i��a&om��A�hk<+�?<@�M~�AU�-��N\tJIZ6�y�-��H0�d��z
�����r�4*�����*\ K�dWԛ��_� ��`v+��i��ԮEU{�Q��dL�뎏�Qv��'`e!(��h�~�R1ѰՂj����c���ה�ʙ=;�Sv!�:b,�K�i&�%[���i���Y�Ѭt�����$�n���[sCE}	�W�$<�!�M�9�e���>ւ^6l��~��,մ�����]�%�>v�/��=�+Q]��GMK���kJ��|���+�������d߰;I%nc� Sfs9<�.̰�^�N ?m昛�!C.�	Ӂ���4�ϗ�7u={O�{�U+y,&��h�9�����?��ÕBX�Y����)SX�h?�ǭ�H�jO�P7���i<2<�A�v,�\��������?�E����'Yy�M��2R�>԰p�]ܥ�����<�vN� v�� -qJj�-n�����@���^5>A�񟤺���禅���N&{s[ks�����ұ�-�|R�2gy` �A@�YL�^}UUlם�O\B'�5sl�;����h)�t�)ri��{h�&H�fU(�#�?��Fβ��a�W�
w �e2{,=�f��m�<��-�hҳm�"-�.�D*I);VΛ�8�Lk��%��n[q�Ww'<S(��\g���	�ew�j��Z��ҥ�����C .�.;�U����\Ih���l���+��ת�\F7BL�����*��,�q���A+|a� ��>BO�;�Q���y�>�"�%t?vTÛЃ���p/�Q"����l�G�*p�S��h�l-�^y\#H�ܾhav(F��_�v势Gs�/*F��:/�d��MX��|�Κ+#zJu�5I�2y�_�c���xY��:"��s&)1]�.�śۏ��R�yu࿑\����X��?�խ4�|���/R����B�E!a�[���¡�#1����k��侢�ܹ��'���^}�|����4?j��)��g�|�@�2H�>H�.�=�����ˢJw�]I&�U~����\'�N�s��J��`7!F{���ฤ�)g�5ϸg߿�#.��x�����,�I_��U�w4�u�/�g���4���mD��2��(�tzT�]�n���̏m�e{pK��Y�a+A}<�ê,�l8]�=zZ_��̟#��_+�u�ċ(����iܶwK�a�|B�����|q���4������߬@��Z��
�:S�P��+!4��n��r�nR�C���)��Ւ\m�wDU��_�w5<&2���/���E"�K�x�u�SSz�I;�7!�ןԍ��,���!z��B�P����6n��\j���BOA��=��xj��aYbX��D߄�m>�2&��*e�����I��á�-��l�ݏ]���碤��2 �XٷlX�$�}���d�����E��k7��g L"s�NP���4Y�lP��݌1 �UXg�D7����x��/k]�j0��Gc�$:��g.%>��Z�+a��[je2���e�>#?�����'���x���FJ��