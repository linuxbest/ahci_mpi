XlxV64EB    3a35     fe0�i	,�2��[t쪓y�0�I�_2��{Mԫ�o׏j�� ���b
�}O�<�n؏d�tX9�����)}�Wɟ%'�Րx��V��77��.Y��0������V i��7�闣���Y	���a2M���!�a�СF5���cP�j��=���ɲ��񜗔�(����=ys�>E6���8��@�E{(8w��E�g�2@۠��B��[?�ݶ���dd�3�2�?�c4�����{I���m;/�Q�BӪ�^Ѷ#B����~f,��׍eM��N��`�:W^�'������ُpu��T���L��\ �#R��9��+�����ة�M5H�Vu�/�_�^b�Sa'���zBT8���^�C���;�An� B�v�&j��~ЗM���r}���+ޤ�Zt�s̔:��Ԃ���$��$��RaR��pm���am��:�H\�j�":)!qx$_V`u�  �wi������Ԡ���ZF�|`aoD�D�:��*�9��x�=_ܹ���w��+T��&���c����!���#�V�-�� 	y�L�dSh����r���п�a"�*��u!��k�z���ȓ��<���10Z'�N2+����7S&���R���pů�o�=�D�@�;��L��O�1ѸU���ɓkI�5��TN�8��pϢu^��(��DR)y�����=�7��6c鲴����(�<4��O�zRF���z?�U��/�k���l�5/L.��/;�adI��;��?�jy���d����i_|A��Wf�a�q	/�Ѩ���h�}"�{;FJ�<с�y������e	�P2ͭs_����Y��3�)Ѝ

(/�-��6N�Rv�a�(^rw��
��X����B~Ž�&C�m���@��Mn;y�Hi�CŇ{Y5��e����6��-C;����1�Ŕ*%���}Rj=Ƚ�����&%Ђ�,|�����07B�!��uA��O=�,
�K
� �����pg�D� �rj��ȋ�-�kO�/s���b?,��~[MU��X`�{<�>v�*�1�y9�y>7:\��Ĝ	R���`�@�=�n���1B�۽��J�C"�?0ֺf]�=����|��u�;�8TT�:�l��*BS\W��C�l
A²j]���]��Fj��ڶ�a<�z >~?�#��'���N��^��㨱	��ݒ���W	]�xf�C~�A!�ƈ��{�#��_�shy��$�H�����.�l�W18����O&�Y���Uz�C�/^B�q��v�u�EO[��g��J5̒A���]#��7���&�j���Q� ���
�G���0cѐ/�L���U�h��(�xV�\�C�@W���s'y��8�mf��ͧyҧ-�p���DRq�$j�,��`���\�������7j�جL����2r�F$����12�$e녪��b�ꛆl^e��n�`Y��g����s:��+O�TٔV��\��5�?ΐB[�ra	6����C��'��]�f ���n�%�AbD��X�g�4�`mX�+xmm<!�9�~*Y|�`�*gf����j/S�\P��J��@��n�2M7�C"�I������~ �2�Z�yM?T�|�w��]Ћz읭�� Љ1?R���lu7(6��/��!R*C;6�^�e��rgC9t�{�[~vw�� )fJw8�0�
�.�2< P���j��!5��|����n���#�P���S4��vW�fz7��K,���	�JΕ�]�|�#�#�ە��N�%LB��������1Z	u�!�1 ��؞g@�F�dY?�컻�)d�tB��h���:�0/"� :�
0�sX�I�!��^�$W���C�a�y8��w�'�s�7(�0}|�>�J�
v��;5��&�P���1�j�h����-�!���D)�α�?[�J=���X+��q6�̫���HYL�3~S�Q�)�,��؏Ş�~2O��`k�V|e)c{#,�{�1ϣ����W=��C�p~v);�1:�Y�R]��nu:��#�����!��JONn3k�.�ЧpI���6=��sd�V��0y�/ׄ���GÎ���H�wn,��)1��oJ��E�	-i��1�P4X�7W�7�)�d�-:aؐ	ۉ�����o���*��̧Z#`����/��-���f���
�n��J���4ڿb��cU>����í��O/q��|F*p߉_���g�<eB��[����,�J߻�[��i�%���o���M����ߠ�ҩ^���g!��K�Ąq�rQ�x�s���U�k��� av`ց�c���!d8����M����t�-4��.&0�ϡYǱ��Q�si!�~&ϾQ��8���1�tkU�E�@�U���>��{�����.�x!(��R���������m=���Z�"/I�X�؝�AF�S�U�\!�tG�
��M��W��7��%�D��7�nB�?��ٍJb>YO��7~e��gj�f�����7h�����ʺ��
7��w߬ ��Lb�TTWjDǭ�
���F�u��Ԧ�{��&h�>��?� ���)k�28���dn�LR�� �\"����o;R!�W�io�t�q�\��n��ɚ��x�n[�Qj�����cg޴��pc�X��s�R���;k�x��bRԻ�Ec[9�pv뵃I�k��$�6O'7��9�?�:�xS=J���wt	�R�W��2�)����cX{�5�m��[�>4 ܾ�h�晒 "z��B�'v���'�i�n��H�x����M@�,@B���Ԇ��9F�H1���1���O� �j�y�&���D� ��p���p���P�\�[����<K�ũ��[���@�2�
���*��<������O�f���Tuv;m ����q��[���n{d} -M�K���E���r��a�s�l>����� a�X�Yu/�"��O(�P�<��Ci�}���$E��B.��/s��4cf�����M%tG[��q���#S6G^�y9�Ȼ���Ȕ��sM�n��}T V[%T)������L�D]�"}��V�d��͍
��T*ǨN�8s�Sʸ�j�l_��a��em��o��dq�қ�����>��w�|�����A���e�Y���^֬s�tЩ4{�;�2,�p�F]�ge tԍ�/��fu��s4��4N�!d���!�S%�a��
��V���݁ݬ�x�b�^�\M�s�9 ��1��4���A���������G"���8���XQ�����t&��"阐�5u��4��g�c�:x�B����MI�iR �(o[J�@(7���i�Ch�	�Yn�Н;�=���W��d�\\[ё�B њ8���U0B�%NИ=��Dx}/C�i%x�Y��F��l��d[,�L�;��NK+MFm�w�c�w
�q(��[sx@W,��rq�B��vR�O46�:vy8֔�K��Q����`}T�":~���>9=X�Zyb�q�>�l�U.�?�9���a�,سNIG���`��'��;4�hsq�tڥ��`9�m���
��-�;�~�o��0�eՑ��^��"]<��x�*���<QR>m'm��B'Dy�R�	M,���CNG��t�ǣ�Lb���~��y����{�ɨ�(���+bbt���.���$��|�b?,�~YXa�q+(2P667��LD
5+ecj ����M�@;d%�%e�m�ܖ%3ql��m2�����Q��������Q��L����l|ȶOSu|�?��M��S{R����4�>���o�9�6�[���Gm�(W�Y���$�Xo(�����kW���D�{�/T�zEyk]����� `PΑNa�f$Ƈ����Ή�N��G{m���n����9��F9�~݅���yP�\ne\�T��?z��/)��6Y���j(r����.��p�FMoWy����/=�(�^G�+v�.��T:G���:9��G���4'�>�}���wCɑ��j�]Y���5������{~ny,L��m�8ҧ