XlxV64EB    40d2    1120�qk������zG?YZ�F��DTM��T�a��K�� �/c'�&Z��kW�|�GV��I"��Ӑ��pUP䚗�l�� �{h�d����d�k����]\�2������-YT���	cx\G�P���E��5��݌WǮ�	�)G+.M�x��rO�z�9�7G*(+�x�>��9�at�r����.�yf̋�Vx@	�f�}�r�FR6�ó���}"@�!�G�ˣ>M[�񘿙N�ҽ�pRY�Y��I%+������wZ�V�va��EL�n�wŒ�ʖ��sуpá���[w��[XY�h��Sc������e�F�� ��Ѩ���n�B�N�5�Q�zcY{�l��tf��6;�>f�
K8�9��>�E��Ƿ�0����ڲ��n9F����<m� ��C�?Z��*��5t!�ʽ2�W_wJ�2ŎZhU�c���h�3��d�b'Jp����;�h.%�	k������kb*__��#��/Cϫl1��T��ߦaw �{���x��Z����p���t���7o{���/��ǹ�즬g%�<8U�ƫr�]����2�v>��M���Eb��[�Ր�U)�܋M"����S>1��۵�3��q�$���v�"���(d
(�VڳZ*5JG��R	؏O�r��
C�&V��[[N��$��U@�Z��+�ңf���TB��@�I[���
-5��?ZteCq�14�ɝJ�DL�Ӹ�av�佦�bc�ڗuh��Փ������z��� �%�Vk-a��eޖ,�HC��\�i�' C�YL(�#��wNpܓU�x`�� a��r�Oc:
���Mc�^ǆ3�Pwk��2S��_ ��40QQ_�N+̇c� �\#�|�Zt���0�pX%���]�0�o�l�t������L���f���ϙB:pH��ٳ���Q��������[�0�+@������ۿ���hݏI���#���$	
�o7jYnՆ������/��n]&�xo��_0�
b����b�&�~3���L�׵��<�i�^t��O�4%��}S�[c���vk�7��ͨ��D�"��.�Tak��H�����yNu������3@g��"��>�m/+�V�l 0���l9�~�T;�nuO;g�ĲNO������%Y&{0s=��'����5���Cjg�i';f*��- � *���b�.��a_e�%aDV�� �̭��U�}�g�����>���$�8���W��A�*�+Q��$���n�1�����A9dօ�	P|�sR_�O�p�Cҫ*t|�)ѿH�;[0=j����F�p�1d�\�2lp��B�X�o��B����Rq�.��P�6���d�c�K���xι�GC0uM�����lE�/鍬���*>��n�O�����m�9�6�mM}���{�=M@5�c��8�uK*g�]�^���_����p�K��|B���00QĠ{��L�׳�f��q�^{��c�q���׹�q�t�H����l�	>Q7��#�3�p1!�C>��rr8�.&wu��Ҏ2���g�,�vQ_R< ^ ���?'j�@Gj�^D��󆸷�oFN���)�#|�)D���OD�v���P՗��z�
������{0}�q7*U�r�J`P���lQ}n�y0B3��$�?�O���d,�ߺ��h�#��e�h�˂��t����9����41V6ss�e{t�%���.u���������^XH6�b�J�!g��%���w���2/��ɳՔ`Z�SqZ������;�9�*��H/�;���)���Kr�K�A��|�/i��|�7bjNXƎDr}�6�Z�F������������z�����F#ĉf��1� ��B�� }�K�fU?I��NO����3�FuMT��+\f�;�v��+��*%Pq�&i�t�xx�44�~7"�a��Ĳ�{����K�Wn����h��Ymz�Xl(�t�I����7�lhG��W�N��Y�$H�`{����NUJ�Jt���c�wxN�hL:O�躌�3Q�@�@�C�7�9���h��R�B(�9l�k��v��
	X�&�%se�-�����o�.˞�cd�H��3`���#^���,ur��;�c�EV&o�Ö��G2�A���wWM���}�yz�*���=i����0�Oo4�qoz�?ZOZ�nT���q���m��U�p"t�$�ϔH]gѧ�,"�5���1E�=4S�W��X����ס/��Y�^�o����#Fn�Z�0y�����ə�p��`��3Mi����b�tn�V.�kG	  �C�`#Q]6��#�~%��xR����-57� \3��\�|Q7��G��An:���T�`��U�Q�"6�f$�7��������������9
t<�E����ʲM+�����D[G��L�>+9����ޠ���qF��$�(�s5Eu�޸��وXxK������y���1j������
��_������VTB%_�3l(�5U��J��LVo���M1^7baI�uf���nn�!�m��r���8B?G�&R�d�������8ۇP��Az�;���"<��Yhe��=K�^�O���r�����n���d��&�^^�T9S��{��0��*�ګ}K�	Zzx�,�75#�� i��]��M�����W !�7$m�>˭%p�u2����P]����wn<.f:�����x�۹�j��������n�ۭ{������͹xeNBP���/�׵�7��j(�ˁ��4Z��>�`I8�h%pI��w���������T�����X���ho��%��Z�1�����{���dn�����L
Т�n�Zسd�==�VۭG��1yVvV;?w�p��Dp���-���������B�N���N{���'#��2վ�q��	����߰V��S�u}y��/,dG���)4`�����D��DN:=
��E�ϩ>�F��g�����[_���!�5��L^Hh( �F�r��W*z�*@�͜vĘ��=Tz��i���.bEM˦ l�v���7�N���U�a�$E�rc��԰��+�c�VS��&�b����ǯ�V%� �ߚԪ.�����b�A:���Ң>�9�%(BҋU~�N=`�C��z�����Bn�z8�K��Ö�쌴$�>9�_�uT��i$�D�g܍�`Ah+�������J��)�85���g���b�������d
�e(�n1�H�}��� �m�G5��Էů[A<Bc۴jA�'��hL� ~��]i+/�ۨ'{�����P%)�V�[Q�K},�[fЊ�9�d���.���4�C8��Q��W�#��2u	���DE�U*ģ��a�Uy�8��7ϤF�&��,xYܫ'}a�eu5��0�/�������Wr�()X�_v�HꄭYG��Y�}�[�_V9����qL�,��Z�����O�r
�e.��3T�
�����X��� Px1ョ$��n}$���Rb�d�u����l��v^�U֧!�l�e����Wڄ�%3~5Uxf�A����*-�eR�5���؁*Q��aQ�j֠m�q�����ٌsl��PS�dLd�mHC7zX��6�P�������J%�C�5[�5e��4��ݞ�'(=K�U2�q�VX����׮���Go��i�ű�^}˸L�,&��jj�29�j
l��+E]R��Q��zO�A�ZKXe"�#@�����9����D������m�T���pm츺1�r�Uz��6���B�
���ٟsH�-�:�{
������W�
m�&K��>��i��(�^�`"X�UU����V�z�?�e0�VQ����BH�_)h"S����D�h�o�Ly>�s ;C�o� D`BD��6�qR�j�G����1�V �F�-
�YE���U9v��Dr\��﷢���m��b�#��R�����3�����>�DT7>7`�v��pub&R���2�,��<v�R^xv��T4SW@݈�U��˅��,�C;M��5/l�5m�`�n=c����M��s"�7� m�o�+�cJN�#�m%�Y�'_h���娄H���+'@!�~�Ȥ[r��o�V�-������1 �rյ!VU��7��p�x�(�}+� �XCf��R�8�x��fZF�Q%^rz��=��"�z\ �Z��ϵ,�M���F\
�b��S|vE�
Z��c�������l��(�d�ҿ,]��1��آ{ذ�Nw��m�-�8��;��e#�՜��9! ��g7�6J��a�n�l�ԩ�󕿊���
7{��amN �S���PO�1J�+�P)���#