XlxV64EB    3bae     f40���yXp��L[�P��zpw��a��T�x�Q�Cqov^h��k�:�S�GS$�]<�޼�eR5侁d���D�/k^��i:J�Q�Mr@N��?Wp	�?���2��yκl9e�� lA�t�j��0�[S�<�e��G�&4M��������eem#8�A� ��I��k}�FF��g��n�5)��:iّ͎(s�B�����<�V^���*o�?(�D�E��Eq�w����!�d�+R(�� c on��߂g�'�4η�B7����~��ts���Tڟ�y�}���i���+j�vFj��{����@�A�}b���q0�3��̘�
L	�ff/�ZSiW]��9�ӓH�
o��.�	�K�6&|�RL,��Lf���na�a	��i��G��������W����?@̐��RR�yq>�r����jΏ��l��6a8'@��	�-��q�h@WU>	������U��f:�R/��G2i���=�3ok���hJT9a�n� �#� ��7���L2��Zפ�Bj�I�[=}���c/�)�zb)��1���jK��6Z�c���%:ٸ��0�s ���+ ^��e��+�U};��zĥ�A�j��I��&2�n	����S˝��'����LʩY�X�����&r)�E�����6�<[.Y���򿊣��j�����ms �B�N���Km�7�i
6/κ'�ʥ� �X���ʯ�V���|���{~L�����'@�iǠd��R���HB��s�"�ު����������,��� zuAՈ4�5졽��K�_�U&�`������B	�O����*����ޏ�#mK�q�NS��;{���:��:(f�*q�L^c�k�
�oҚ�~A�<��L�$�1�W������xo ����*����Z�IEz���H�GCIkRP$�4'�}xZ�q�qc��\ ���D1���+���fk�:�R��#ꂸ�=<�Dx8�0H$Y�'���H�y�2�)���P����� p���c]jv����g8T�243[08#v(s�V���-���g�\&兟ظ�͐pT�A{����5�u0���3�-t����Oe�c��B��j�(��K$��}_��'�d$9Xs�!�:H��/�٪���i���|w�}�����8;�y�6)Sβ��	R��2�u�ע�����m�g����:ޭ�wp|3�SY/�a���Jc�&�K܈�hJ��e�M�c[AeIh�m(��qT%>?��`�D�:�M����O�\_~�W�|`3��ݔ�C�[ق�����*lXS ����,Τ���h�����ޢR@��^k���zh/�^zP�|/m�F#��2��;��4�M�T��\b>��&���@������$Vs	�Y�W�H<�M������G��z�Я����9�M��#���u��!���䓩�n�����nm�iD{��`)�ڬ��`��+#�������k�|�Ir^��,z�S�P�����zī�jH�ƪ&�&E��oȐ��������=_�X�P#��:b��V ��x���t�)�P�(D~bhf�P�%	�K�\��І��d���hP�6�'��4ԀKk��7��ꚋ<�d�ȏz�-+���o"�%<G8�қ�\��9�c��Q ���W�Lp�X�Dd\?[g�U��~�ѩ�z�Z+��>�O���=Q0��{�i'RN���L*^`c'��{��a�d%O����ϡ��ރ�}id{�[�K��Li"U������˛�E�p�@>�gOC������O΅rdhZ4ૠ��e�;&K�H͵�����B��K�y=��������������}����X#����g�Q'��Ds��z}�'�IFЙ+f�Bh�l���daE���8zd����

�׀��SӚ��"�����8O��1{cK����R�|Kӥ�yC����De#�z\�a�d��U���$/�-��I�����$0C2�ߩ8T �|F_}���w���]�5��-��'�i��[|2X���������f�g7���(=�Y�����j`%Nԓ�p]���f���]����w ��L'{��ݛ*��4��݃���x�+ ����������=�L�#M�.�� ��v�HJٿ�h��k����Z�?^���oGeE/���{�1��|�*j$��"^͠ܛ��@��P>l�@�N����ƛ(9l�4��Z]f++�/TJ�ӿx��pj�6��b #�wBҕ1�D���jm���(�f�F�m�d���-1��G�f��N�Y�x3׹k��(��Pרڗg�Om'��90n�V�;� ��.znvsBxu��q�� �p�k�} cM���mG����VB�f�y=V&���
��D�����G�j��H��oo{-,RH�H�����XKƻD����EoG;]�φ%�1��nbv�h ������SI3Oz	�t'�qC`	�V��(���\ux���&cIiI3�Y��e��D_Ż���!���I��/��HwL�]^~d6��7YT�գ�5�9"��5Jv<&XP�z��Mr�+�8���Q�5����0\&-�ɾ�lCD��x��k�ۑ���?/���k��2�V&NoB���w(�5�T���4�Z*�_	Y����miTy�o֍p��x�#G�Uf��9ڡWS��ꅦĿ]BŚ5Xg�O�����B`�0���t�'�����5����>��AYf��_7EAW��P�=X{+�R9y�i�*S��$cOu�Va��al}p�r=��"O�(��v�HW��}vRp:���芉��٨��o4@��[��ۮY�w�f���K�������|KY��l��~�}W<�U�-�b��H�(
2!8�E�e�!�Zt؆�� ���#Ō�5�&��k^7g�Vpð����l���2�.5�I_(YU�SP4��Nޢ���п�ϧ��6lʆѓ�=�����&��?3[x`_�BX'����%5����7�0��֦qozY���٠&��x��q��ϱ�l�ҭܕ-�Xm�����Q�)Y��Φ@�]��@�\����=�>���m ����OC�"�A;�����ȍ�`ǹ����ܼډ�X �,K&k����Uo7}�ɰ������M�������T�s��s��HL�c��D��D�6�yc��T�_7�*d�u��
�׋��K2���pp{���^^�X5��t�>H�������忍x��ަ�$9:Փ�M���Xr�8�a�*� 
oc�̭������*V_ğS� >~h�}��1�k{�����ו��!*̓2���?��u�.��iM���y���wY�s�I9��0�om��b�k�WM��Lw��� ��)�nC7�v_�
�3�d�s%�+�
XmC����jEvYSd�M�#��4+i���N��z��)����~ bh��k�
���꼗!��q�%���Ӷ.�_M������V���N͐����VF������DϤ��@v�d��s��|WA=1�쪪{���O�`ڎ,�\�H���k�U������3j��\�>c�-�ǖAF��[��Ey�@�<�� ��J���Ó�\h�R �;B�5�������ۻȔ5X�0�c�vp�Z|����M�(M �]H�@C��&�%A��}��oS���h�;k�Hu�&C�f��̻�1ڠ #�?��<�t�$ǜr��y��?:&�d g��W頉��g�� ���l�]���VekJIʦ	��3?T��#����F
ܶP	چ��U�;��T�o���6��0q����n�f�����্��_�L��v!��0��K�V���.A6��c�K�f�