XlxV64EB    fa00    2f70i�d�@��<K9�^�w���
0YS�A��C�?O����%�5�K������bxF	�EU{3�vl
V� �+��_��'&�zQ�����y�ŵ���5�TI컸�z��6Q�#20�R��x�?���ٸ��� ���"�����B|��Z��"�s����>EY�I�8U�pd��� �Kzm�YYP�6��(b{�N�K�-w<�ys�,��:E=τ�ʯ���Co�s�,M[V��c}W.�D���Y��)�1׹?1ke�x������e�Q���v6D=P�9b	+Dh�M�Oi.B���� �����ίc��*H�����}w�ւ@p�����M�_x�?�'@��e�	_��֢�G��%�]��Ʉ�KO>
U>�Yf�e�<�`,��Z���d��0�M�!j,�,.��Q���ᕷ����)o�����o1���o�O�hL�My�}-�� :	Q䐄��w��/��Ń1�v#F�~ �ɯ�2�j�j|ڱ�vj��t� �ia�A���ޖ�3���+L^��B�]����?��F(�X��	.6���bL��8O��]���<���缐�$�(�'1&����dM�|�:�#�¾tƞ5�����f�@�uH�ksu��$���T����6b�^�L���&���E�l�|��O"�OCt�kЧr���E؎���0�ݦ��k���7�Үi��\s����9�����������+6$�����*~<n��v��+��
L�"�3���PO�Ő��t<XI�����bS⽌�@i]�/���p�d�=ǝ�0 [���;T����i�J�tc���U���M���0���Y�9'�H�0_Q�Ì-4�L�H{�X�]��C��+�_?�ʋ)a&$AlU�	�r]J^
��T��� ����F�6�~oj:Fn�%�m�T2X�'U�yis).�paHV�:�z�͐ז�(Yf�K!:e�l�����[�B^�i�kH�a�=���n��R����?����vz��@�#���"|M�8���['�ܭʔ���Z#�/��-��c�����9��>O���X�j˟^�n�u��G���j
�:��#{TW3('6�W�Y_d�z�gN�� �T,?`L��Eu��EV��hs�%���~r�m���>����Ǜ$)/"��IÏ	��= �����F�M���1|�����/��@��x�v-����wس�([��jDޞ8�ߩTp�N��t�Uэ\F-�[5�&y>or4G����B;���X��Srę�n�,:����L�7����O��iP�����"�2�Ϙ��I��7�?%ʯW�б�B���<X*.5��g�P��\C�5��7�I���<VW,h��w�,�1��*�P�q����$��PS=��?��>�Z�y�U�����)d*���HO����O`�����F��%M�k�Ra�^��U�dA�RJk�u�!7���$=�d���C_��4�ՅX�Zw�;�):�e��Ŋk:ػc�;�*k�Fe~)G'���'��A��ME롊���h���@o��kF4�0�U���Uq �'y##�^R"+��l�� ���-�c�{�&�����	j�27���Ԙ?�/)�*�k����D{��ho�{	ۘ�LL`{G8>=^e>��
G�?U����M����w��}�z]n�?+��@7yI�����f6��|=��g���1�$�®�w�4�N��\����>{g��J��#k(H˃���q��(=��!���&S�G;,���Њ��R���#Lv,��02��@~��к�f�3��X�@��QP��E:N�q"�p�i�a��.@�T�\ A�����	����V��'NC8-qӨ�xt����=t?
�@��=��c{%8%L�w�;�����f�j!�a1T,cbF�9��t�Ǒ�~rS�+�����xE5�6�i���iCT\����ڛ���R>L�<���T�F���r�u���]���	j�J]^"=�x���ܣ�&�Sae�J�94�ڲ���=>�QΎ0�E0�w��"�6
~%ߢ���{��p�z��H�yMͼj��m�1��T��VN]�Qn�R��{F[��b�3����H�];��W:�3�OI�9(�p]\�H�5'������;�kQ�ϋۃe�֏W�CE�G�X��$��s�BO�\˻���[#EzHa�~6e��Kʧ��_WۇK�L���s��-iSU���������B7�@��4�2�C�eM�Im�cȇν.+�E�y�?�Z�I�и�aA�==�Ww�	��Zo}��
��Nͺ����h�\��t#�Z��,�L�����#̄R/�`ǈ[�ƺx� �Fi41�/ ���"��SnӃ}E�.3m��Gx,#�y�b��C׎lSΦlu�y��qE��0�(�.��G��}7�Pz�uVGy���n�;E_������9|/G�+�IT���n�8bP+lb dDS��N�W��vE�˶۞5kx�L��h��V��-!�F�0g�U��8O2v�q��,�5h,O��vF1'�3_/e����נI�T��W8��
v�������v�v7^�LD.E�$sb��tH4�V>6����Qh�I^���D�J�l��z���,*�+Ҵ��{-��w"K�'K�l�� uIDї���YÕ���� ��#k�� �B��3�C�v�{1�ሱY,E���I��u�r�xWYB{��A�B)k�|��2Rc�X���P�6zl]_��>'=ҙH�k����K4�d��|2��<j�d�u�z�y�,՗��N^�I�����z�E��x�C$=��B}�ƄhnBN}k��B)z�+��͞����L�]�JTeý=C᜖��:�SL���qD��p�(wC�w�{��/,�d'}K]��TN���~Q99�Ä��<b�my��x�T��Ĩm�(�m�j�\jC�`�s	4�*�~�j�J�>��07y�òze�Q��`���}���M��5������B0~pFԄ�������f�u��fޣ���NZ�`��["#�h�V�!���K��G�o
J��&�+&t�:	&Hp)��'�E�����io~otrV��;����uI��ޡ�G�l�1]��S��so*�Y� E�ۑ�֍QIH��z�K�C�埦>�<6C�:<xx�{?��N��fH�",(���3��|�%��5�S���}z{��]�>m�.�O��c��=钟�� u��h\��ʁ/��[��0�Ic{^��d*���y�}w���.�>��ehnM	���M����d[������u��'�/�SW������8Mfm�����L�sIU�{�Y1�����2�C�zY�塒$�@:��P��;C������(S���"\ܷ:� `�pPۭ���U��n����j>���쀅��\���غ:%"��@e��-Ely!G����>�S�{��o�?���R:xǡ�5��!N�?���a@��[b�4q����?�9�?�{f���)���uj_�k2 ��I�Ѥ�i(z���P�EA���K�P$�����v�˸4Ě&�qJ�`�Ο�	��#��!�����0
V�?J��h���{tØv�3�R���@4ݯ����h�����+�)Ш�"{q �HQ�(���$p�1��!HjH��s!���n��FQf�� ��e�o���L�tW�.�})��d���H�Jd[�|�}$?���������W@�����=���7�������͟��2��;)9�[~O?���=I�N^�f�6��ԛt��H^6d2_N@���EA�@�1�,iщ#��˧41���j��bM!���c�%uh*G�Q�O���
�Q����z�W����a�"���ln�";G	I�jI�f�#����-����������$+=�P����R��fzu�ֈ�Ѓ+,Drz�"]6�P��do�`��D�!v��j[JK	�z�T$�yb��c,vw��&;	��}%�	n?�.߾�573��F�5����d2��M}�'3�~�
]�46�V�M�����7���;��Ѥ��C}�b@)DB%��N\��Q��Y����1���)ZY��b�.֦�W��/�
:�^����Ï���!�"�m�k��@��GFO�Ԛ+�ˌ�9N��p�_e9����,���(b�����L*��!����0 �LO����k@A=N��G\^ �lv���xb�H�L�K�-V�����W�D;x(��U�c�<����8+�&�i��3��3)$��?"�a*�� ����+�wJ@�v!b=���
d�l
�Qm�wHʘ�n��hSZЯ_`�G�L0�
K�"I�!�'�q(_�?��Lx�uK���ನR-M�=HR�s���(��ݠ��6�6<"�Ȣ[��� B+Hf�=���n#�z��($-��������}�ʻ����M���(+�HyXhX����]�p/>j���5 ��D'���;a���O��0(�������C�!2> {��H���d�d�
�c��y?)^�/������;��y�w��L�]f����S��b ��o	�>�;��l��h�ZQQu�*\��y�c�s�*�e[\�	��S@Vw�7Bi�
�����È �YI8[���_�H�8��������@/��u#y
�b�O��r^��׏�Bg�4��RK���7�U���[?�ZR��;���X3Gޏ��6Дc���~��>f�#�=B%3�eW�/-at{Y���GzvI�0Z���y��6E��' �R'U6BEye2��k�-.�kp�g����`W�87��9�l.#���d`�����ְXx`IthLh��ka���D�w�
�bhHН��r��*ї^�d.�qM�Ro�ۤ�e���8�AH
)�=�#pLɲ�"0I��:G�<7��R�%;����J��I1?��:�B��S��_�Wb�H��T�SYr)PԆB��&�0�C�J$��H��O��P����:1҈�%�հ�����)�{�}M0���G����*��{�ݱT!pb��k 1�a�D��}���a�GL�w�O�$�޿�  <Q��:E�6Q���8�d��,Z��w�j�&QUP��3�K��� A��ղ/��:�d�]"~+ھ��O�#[�W��OgH
�=T³=����aM�ByD��q5��}R���aIhhSo����Y���G�lDYA򢱿�@��|x\�\���,�8�����h}&���1�K(m���JΙ�����ad�'M`K��&=h��v�I9�.���aU��6]�>U�����"�`-KF؉Z�e����V��Ų�`p�V#��=Fç�3m�7��t���	��Da)/�Ӷ'Ej�7s����n�����k0�����zV\&��@)ζ~��t���3�E�1S�֜0���J$��!X5����9&^س��ڡ1S�I��X�;{�t��4�*¢� p�bJ���}�|������Q���]��4���� 86�7mٕ-^l��I@��ò��7��i����W��;R���U�!�ioZ�������g^�U���������/�Y�M,��q��H����/�tQ�`61�p?Ff}�ۓ��Kj���2���̒"͡9���ۿ��,�$��Ð�zBs��@���`��ٳd�Z\���aPi��i:d[=ݹ�+�S��_�3�a_�
�uȍ �bj|���(n�y�m�e���������>څ�9Xll�K�s6�R.������*�y�+@zm��!I*�):�7^gM��hܩo>��Vvs��O.#zG@�����>��M���Hda̜ʻ������d4��.p"�!6[� ��E��e6�e�2&Ϥ�1g:8q�g%RSl"�Nl�����R����]7��SV��N>ٽ�Da&=�s���H��o��K�+6^�0��
�By��K/6�OV��T�����Ҋ�Z �P�����5�J����ˇ�T�!��\5�T/�{$p!#���##�w;��M����:ф�M�ڴ����t�d<��ITD��	��%	�x8��;�@��M^K�*����2C�����츁]��5%|g�^�������^�!d���	�`ʜ�aV��	)�o�H���6����}E��&L~�6q���S��+���ӮvҸ�t}�ǔ�߶$Ze����{0���M�9��v��"JE~�"�S�&;������g��8��~���-�k�����yD�b5������9�ж*tϰ�p�{+�@X�^�s�����f�
s��A-��.>q
����*)����C�ߤ����3�K;�"jlƸ�F䌮4�EZ��9	�Z��w*;��m�n�%������I�ɵ@!�Oա��*�A���7��_V�X�]�K�B[��|)L�v�c�U�,�?���c�'E�͕6|���j�ɍ4K�OkW"��cI�SN�F�T
"��L�wx�x	ݫ��@���qHQ}��n������DSp&���2�/UP��A�����`X�����Yٰ*��5]z6}��^��Ŷ6%9�*�/+h�J�n�4��7ޠC- �z��Ce���i�P=d�^[,��$�`
@��ǅ�-*&�~C�<���.3�-*����˵�0�H�y�Jf��pg��=͊�M�,r���I|���iojz�G)|ksa�+@q쿷�����He���d�����V$���i��Ñ�����$����#'�RZ��f|�x��vl7?@�t�V��Ⱥnd���&-\�k���E���⤅_4;� ��S�J<���0ߎ��"Yk
7���6~(�zԨ^��@s=*�^�#]�u��bC*$5�N@���pOYIGº�>�B�$л���qSn ��ME
�[�"���B,7Ch�,P��1t�8�"Q{���>Hi�Zi���V�+�'o���'���P�9^�ܪ��`7Э���B@�m�c�Q��([�F����!N�JPت�2��wyEQ�ח��~A& �>u�g�+zi�X�fI���ڋ%�1�MG9�}l����_����=�Z�������is�+�|H�|o��r�N!�T+�����g3<` ��3%�{��,^�F�x�_%7�z�	ᡱ�J���JJ����8+cy�U��6`z&@�y�+�&�ˉD�,�*��kL��°-V�����U�Ӆ�X�$V	&����ֽZ�v�~�q�D���G/�}�'��"8��(������Dk�JU�c��	p��nA�P6<Lp�!�ߝ�
���!�NA�����mkCדDh�x<�eMlx�
���d�ݏ��+N�0���#�Q��/�4�������˪ݽW���up-��*�� 7=����4�����[H�e?�v���5����U�w��
� ��e�cw�"�۳���*����KO@�0-]�O0`�7^;m��|Q���Q�CȖ�
q���qo�s�nJ�A�Θa��#-�����@a��5���d ����\�$�݅�k�k����me ��8�v� ���7��������8.Vn�R2�pVPa^$]��S��[ₐ�(�fi��߷��"G��`S[0Z�Afx��?�f̬���˂�E#a*ƥ��-9���Ӈ�k �(5����W��'��,P�رV"F�7��[����¹y�/�d�k@l�B����J�M��^ǀa.�a������ݛ/�M��i�jH?>腐\����f�zT��Q��U�
�o��k*~+IJ�m��]�{�Ӿ�>�u=X,AԳWi P'.���b�FSor�b���8t�+]?�]��F�Q4"'�oo8,�s�&���ۛ�wI�T�ڪ3��:���i�ӫ���6�3z������!�ۭ���e��A1���K�L��X����gx6q�s�ۍ���~�8	��+�#��R1�%�N�`׮�QL�:���@0��m�Ǯtwt���Z,2uo+���9��´ق�=���� ����6�}X,����"VJ�S���y���G�G	��q�t�3$���Ʊ1��:x%�������!���m���\�_Bvk�ٙ����w=�D����2FU��M���XX���c�E��-C��j�i
�Xn�q3�p��֨9�����u��*���K�{��ȭYUj�`�&V�a('(�2_wì?��-�!��M�U�cP�+���%ȏK�R�}�f��[;�` c���}=��!NE%���	/�l�#��E����
�~9[M�Ңz��6�
p��1�xِ����`�G�mK1��+�܍�OiZ
ȸt"HuN�D:G� (C�g���^����'�&o�VM������s{T�HB����-���Ka2�p���6�E�Ѓ���@��Oy�.K����D�
o1�x��TmE��ox��!�Xv;� o���2���o���凯$�hv�=O�_��;�s@��.�^8^Ɉ9G�@+�c���Vwl}\����C_��d�׀Ҕ@G@ �81����k9l�D�yύg���q�r#�k�z���G����ǘ�P=@ᲸŸ�R�-�#�3��o����3�F����)�~Li2��)i��R�w��^��C1=�ZjA��b�V�/��B�̠��3)��~3���l<�� ?3ϙܢak��g��
�K�����-# kg8a�L	*����.�Ro�w[���M=D5@H�)nb�!�E���юX�K[�c�zv�^�4�d_�$�kq��&,��X�b��3��kY�h�FL%gg\3?����O-Xh���׍�n�\��:��n���Л�e�=9/l&���W#��wH�)"��s�q�ښ��,8�ѥ>{>�T��r��TVE1�(��X��s.�����1�iޣ=��Mu}�2ggC/�$X�6q*]�kQ��#&��ܐ.旱%Ŗ)Ƿ �ף:�C��v���7ZQkd5?ft���g�oh䶬�r�)���~�_��75\ )+ �KȜT=t�KK6�����f�cPb��m���iTwΊ�<mZ�k%i�ǹ�p�A��bx����}j��^��˽��]��2	�&������LϡM�!`1x�ӧ���9T]ٍ\��pNAE5�$��0��!_� �T-�C��@ٍ�n��.Fן��K�˔�@ՈSh��v�������Z��$���N�"'í76�d�W`��W*m=�d�}<R�\!M��~i�p�M�'�وҾ�u���Sl�4�\}y�I�7�r�Ybǖ1��6�N�k�C�7f���\�n*��͕`U�&{n��^B6�e�f$�g���!�
xr�x"���.�#AE��$��ő�%��M!(��Ӎ�3�3�U5+l/����CcW�(J�6e���e���p���&��x�Ԃύ��.j��@�,�+���8��m��R9�B�`B�oz�����kY5D���������I�J��2����)UyoZwA2�X�]�8D�ݓ�!�P�k}֘쟨�뙪T:^\^��l�)�	9Z�����1�K��;��IFu�#\��K�����xv�Q�F$��b?`�҅�馜1���A3���L*���]�� ��G�x)oy��.7a��f�9�B��(��?��.�H����%��*�HP���n�sY���ve�^��=�"��b;� �B� ��W��2���
X���ʚ���'���ٚ53����ʛI�s�@eE�ǥ�Cj"I4��Go��GLk0����W�������I�|�ɖ|��^��`oO��*Yl�6��]��ܷ}�]@���7
Jh���Q8S�pJT[�$c���	:�j=�:r�&���O�$ǐI�u�x�]���C	E�oW�{���Q�A�`g#�*\���b�xf��	\��6)��b9Wד���kAJw���`��]���H>����ݠ�P��W���x��A�R�	#@�k�Z�":ڈ��b[�d�/%E�I����[_kwI*���	�lS�ܪ��/	'�+�-�����Z�\����ox��I8�rq�^�]��[އ<;L�Q��(o��� ��_��<�b��S����l���F2��C6J 肖[�{�$� x3��.R��ݪ/�� ZGIrA�̘��`��r��y���?��
�,u��9�d6�<#�s�B�e�.;��.�<��/� ��C��YsD9�j��k}�X2%���S��"�p�%6�؏���M�M���M\Q��:�/�.��������{��[���+�=���~?�g?+�a��G�p���`�ڍA	y������}�J!�C2;��`�"�2њ+|�Sa�t/�E����iUӢtpO�/<���pTql'!p5%�u�3�ψ�� ho�÷�x�EF,5{z��ln)�$�V�c�	�x�R����dE��jv]��:���qE�:��sö�TG���V��;�]RPU��y���3y��Wu�ꏄ���d��_/(��`��u�E��_Hc���.���>��2�>zA~��ոD�fv�	f���u��Uf�`�+Ϊ	��!���wgC��1P�w�Q6�\n5.�C�蕦2��]g��h�R8�N���ZC���P�m��ֿ$�G������߃�WM���):�?s�-fI]�>�	YY��O;�"�����((7E��0t���o>�F���� sI慫�m_dꊵ�r~��cڪ+��Z)�kZ��~++JA5�))�4��d5��y���j�w�
��V��}I%ƀ&?����}�|�K��B�X�L�K(�X?��Ƴ�$5�(O�R�jcJ�,�`��4C�lQsxq/���V����4�M#FX.�5I0��ʿI�b��=�Ok&�,�|u���2��Q��Y����������U&�Q�I3q+*�-j���h�JK�ֳ9��?�n�cXej6)�����ëC���D;R�,�����=]�n��6X��.M�e�� a�$�Gt�0���Ѳ2�H]���%|�@v�W�rKF.���ɺ������< �~�`7�lF�G�]dt���u!�B�0�����(��ΰU�f�$�ti�uR����\hu��:4w��/�P�o
������w�]I�Q�ျMSGIa 2�m��D�9�_I��֬�1���.q0��3����判�B� 9A*�M�_�b*%��8����=�Wi������S;�D��_��m�Ѐ�41�($�}l !���݅�@�={��u����c_�Ә�	��i;c9Ѹ�_�0dI!o��Mݦ53�W��Ү����z+�_P���S���ϒ²3#E�%I����~/�S���C7C̏'��.�P��PH��W��A"��s����C�m��^��1��V2 �Q���cI����d��&��dgA�j�oa�L���4t6|L�6Nۇ��2S9��W��p[BgLq��6#Q$1|&��@�����?V�����s�L�q������P	0�>�&>M^(�q�i��Yw�W��M����DQ�y��{Ĩ6:bv��¿�
�I��9ژ��b4��H��O���2F�|��3�V�_o}��hiE0���%��%՝��S�&U�7-6����ޟn3s��֬������_�Y�����z�H{�)�"�;e�jet�����ę�����qi�ҳ�~��+��
Y;��*�*��g~�G�A8�Wڙ{�G���E���c0-s'5��MD��������5S��mA��U���,T�o�wn�?� ����3 i,��wg�(�02�Np5)���p�II��(�Z���0�'��[�}��{*�%�Q^�`}�Y&"��Br����'���2*Y���} ;� ��2���X(�*�~�_�G3���k ;���cjrĵ��{��SC��yDML��M��<7����Y��ۆ��o�1�Y�8ClYiXlxV64EB    7a9e    18e0�7�`gwEXe�\������X��E���iT��p�8���h�e��v�uC�#%��F�$~B���IA�����i������:=��d5��g�����h�P��"w�ak�(��燙����gh��2����b��Ac8����|�a%fX̉ ²�4~�L�Y��`L�"GBx�$v>Iϟ	Rb�Klhv� ��es)r��%���m��!�]P����2��)�y�,2A<U������R�n
.G��;�]p��&��3Ay��(�{x�Q �0�N�t>���%1�!�;X�X�?}���ǋL�ꮩ��˾6�/� B��Z��D�N�^�#����_}O���"L�[�7���[��%�Nރ����v�|��0)�.�H�neIט�eѶ��Ծ�u���-�|+ܼɜ.l	^$��gBg���ZX����C��!�;Ky��gz܌�)̗P�~�=_]nb"�h�W���S2�ss��?>�D�Vo,k�j�}]
$�^�ݓ�1X[�ܽ���.�z�(��f����(F7�nՊ�n�F��Q��O��]�<E�D1�.2K��c�a��gH�u�ۘ��3����t2h ��Ld�!f�{A�5������3��`@3��)�9ڈ<ׂ��K J��b��[�3say��K!{�㇂�	�w����Z|�!J3a޾�I$�Ƚ�7�ɻ|��Z��Z����x. »�w���'X�sԣ�cG��T�S:�P�����֪�j2+��~�I��0L<TqK��+߷����Uˌ�K퍜:�3}6>��T.��<9݋[)	��k?,����t�� Y��^�p8~�iZq�Y���?�`]���yG%J�Ӯ��(�Ǻf���I�QѤƦ�����@���S~eH�����A?��*%g�RyOH��Q�΋��e� �?K�Ҩ.��D��uךkw�c_"��iC&=��h�;lep��}X����,6K�#?q���g�(�ކ�+`�);27��������t�172�YHs�"@q��i�D���������	���o36@�h���/*ȍ�JӃ��Wj-�a�"7��_���S es�w�Hv^d8c�������8x��==B�4��j�S]�wk������I#L:*ւ�:�Z���"�26C���Җ�7]�e=(�
U����4�>>P��Q7{^�U��.
��yT]�(۟b�=�JA �%�hu�L� ,򄥿�b��pmv���d`͘��$�g�v�m&��}�V,#�C�#;"r�x�T��D��30Ky�8,�ϵi�B��I���?��l�]�k��`>��V������"��}��/�k�?�5���.	�7���P�m����ĸ͜��f�2P�*$���5K�2��F8^��,���75���H����)J7����@0�A���H�el#^ݨ�ۯ�j�"�V��l�B�	��+�J���q��¨Zl�JZcC�� i���s�NƺЫ|��N@�}v���a��=�:�� l�& lg�ʵ��O� ���>����������7�b|��"#�,SuWS5��&O�ϧ0�>�Vq�.M�m`���~�-��=�M9�,W(%�C*7T�R��w�	�^m�t�(�F9
��|�T�Q��>G�m��,�K$cR�=�5�2��?���⋯H��Ъ�%�˶��Bz涽"��S��U��u0�h%���Oy"�#A�k.42d8�w<L�6��(u h����.�@L��+��&m��qn��U�l�&��>zC��?�$*��E�������3���~�� 6܆������T�L!��yc��&�c�¿r�8�M�t�ȃc�fܳ������U�Je�NG8��y��z^���Q�p��Z���ߘ�E��Ǜ�=7�:]�ܮ#��Պ�:�V�H����
W}�q,�f���j;��~'�鬐ǬLF-T�$�t�r�j��#���.�Ia7�.�<�'��������{ ?�]̟�Y�r�K>XY���P�8�ƾS��P]#q�\���Ty�;P8w/�'?�ƹ����z��K̵"�v#�����r�l��Y"|�m? �t`Z��+����x���ߑga���0��������Aޜ9��M�D��h��LP� ��q�M�$lzg*mK������>�M ^�[5�Y�Fu �Kň��g� ù/��M�.���B�[	&�'i}j���Ku.��Rv��#Q��6[�xJ�F~�c��	3`g��[b�,���Mz�^E߳��P>�I��7�?\�\O��l\?� ��9 �=��k��B�z�q5�@;��|�Za�A:sA��D&���1x��\�q��ܬC�N���?q�Z���E��E�Ȋ)�a��Y�w�C��'�m�����;�d�g���|R�hՁ�9�^	����H��Xf��j���h`гx����� xBFw(J쥇��o�Jp�H֔`)�m����3��2�DIm�8�<�Y����?,� �?��:�s�%G<�V��*
��l:̲���R�N|��rA��ǖ���'~�l*���i^U $�@���dK5��S� ��?E���L��`��"J4M�ժ�e�֐�y��wd3�K�u4�rp�_UP���تbޒ���(�ʱ��������$asQ�|��Ŀ�X.����
��lF���Y�<��;�t��40�D��|��sĖ�V�E�TO)x雯#�o�����ak���I�_�Ŋ��P�b���+�l�|���&�� F�dW軀j��l{bN��B��e�2$�u��=FWl��*	�Ʀ���7��	59���}DQ��"�;)0.;_0{ۃ%(d��]��r��Z�}of��];:=D�{WP� $��Գ -M��D���"�2�i�EIO����I�AĎ@<��H�s�$K�p%��Ӡ��ڷR)[fk��T;�V��K����y�i�Q�=Z�]��<��{"��%v�w1�T����!F�Z�q��[�V�ٮ�7R��E�H�Xqť���������{nq�c���K��X�e�`��Q�uJX�;o��񥉔Ս���?3:Z݆�m��eyp���7��R��;Ph�@�&s��I�+S|��<S�_*�H�4J!?hߣts,0����W�U_��
G�S���xD��_5���6��[��bR�nz����1P��d�l�D�4����H������}��z�7�R������K1]7���b�L�
�q���s�>��ea����l'��6����I�6��ˠN�i��=N��+��b�
O0��v��M�#2C���[Д?t��	lG?Aȍ�X�)O_0��&�%F�I�;�����4VV�x�׷F�ʦ�̥�W��Z�3�����LZA�'+q=k��q�X��\Tܒ��@�W�}8�/�(�߄��~��:��c+ *�I�?�DP{�P�l�B`к+*�����������6.��w�5J�@��x�������@#d���e��&��xJ�9�+#�:'�ݧ?����(,��1N�uA�l��т����?���>e��P

��THE�%��" ^s�b�FD���O�pqRG{/<J6'��ʍ��4���ͬ�ǥII�e{�S���%Rr���;_I�73��L�6)o0�m��L#�L��b�g��^�T��B�� JvЋ�	UV
�FX`���0���g]��r��Fg�1�N�xaw�g��KQ��W��k.x	���I��6'ڝ�����J�gֲ�||k��JhO4�C���s~��X��$JC�'9n��n΢wX|4z��<KՄ{�CSO�Z��)_��g�~H�ݩ�ѰI���;gq�D�����簷���,����P��{�o��։<0p�`��zL�v/��K>���O�km�߂���w*Z�W�w�(k��|j�d�L�TX'tJא�s!u��m�[�����07o���fV���_��Di�o	
�K���d�+�x���YƦZl�3���e��#�Ᏼ!|�3|^��A�m��V�,Z�Õk�c��p'��4��W���%��)��8ԗ�?�H�3�?|�۴IL9R���Z�7T�m3 n���6[�[q��?C��<BW��U������An,��5�e��=^��N�v�ʒ�׽X ��Vg�����U�6D��2T4�I��4@^�A����|#�GG=e!�E����h������qh6���;�^PGԴ}t�):�/���aMa!z<� ��������1�E���N����R'oYwPxu�+������x1��s�M@@2DC�7��'_"��W+��wI����oF>�ܓ�j�+�
�<��Z 8ɹ���s�Y*�p"��q�3���݈��:����8�KD��(3��rݑ�hJ;�E�4�Zʽ��Mˎ&�$0��Z����DM��3wg�>Ϯ���2!f�j6v���Z[10f�}�L���X:��"\b�8��g����oB�&`�53���Tz`���+Z!�k�:�pfJ�[��c�4^��6�.$�8��S �v�,|��P�4���[_S�yCAhF��!�{�M�� b�o/��$�N�̼"��L$ڢ̙`���f��ȝ~�m3�Rӛ�L��?b�����҅�� �]�⫻ʠ_T��6�G��.��`��d�@С�N��	��
�ޞ�.|S��<������q�`7u���,bJ#��p�O���@q�#����<԰�X?�/zU�5���*����M����#9J.7��{����J�$���n��<��z���;:�]l�J�©tn�0������j!�3��0������Kߊt��#u�i:!�������^޳��7�l�L��g�U�&��oV��x�K�ŧe�!��v�7�JR('���f����9�-�/RH�osV:PI�m���DkoiYxA^䰤�
����XL��C���Eߺp����)�0����ZH�د��MY� g���h&H���
����a���dz����+�:fϜ�)v�$�����!(l�%�A�e�}�B\�T5�n0ߏcï("iS@e3�9��Z�{��۵ �	PX�-��E�G�ׂ�鲬|�Q���$��Q�����������%�$1JU�[���R�%D������mH��r�������Ѕ��RK)���4��Y>�쨡�mZ�T�va��zF�c�]GC!�EK07�����8�Ў��Q��rk�7{���N��kr���>�"m�|�ɘm����P����3�,��ˆ�=�ƯV`��~1�덖M��i��^^��|{ �&�z6X��o}ޒ]��FC����Q�*���&Ut߹�ڻ(wW�|��@���/CO��g���{���� ���7.>/(��BQ�!��tV��36������n�l8|U�F���� '��,7N�Ja淟�つ������˯#���;�����%E7�Y ���\7��#�?P�^��/��!�J߹��%�"��z�������g5��A��U���?�(��񲜓I*/e&��4�C�
������j�#$�s� �5Xn�C4��#�ؠP)�0��}�as���9�v���j�Sxƨط��o���9X�\����G�BXG�S�]�|r ��ɤ�:20�Qu�@v;��C���$3�h�?s�q�",�ǝ�E@��<�g��OU��Y�6'��Q�aLgD7}`:#�_lj�_d~��,>?��(�Jܱ���y�Ҡ!CbzYh�'@Q5��<��,L&�Fb^p���v2���Hwb��z�<�`2M�a�E=1;��+�߮a�u�'��1BX!�ܢ5�"Y�A�H�i�K�3��Y�w�r­��E�n�hN9���J

�
���.)��盁o�7�z	TR/� ��ڎmP�����!7��(�� �-09a����eJ�	����K�1JSÙ�z_Q�z**�˽�`|^qwe����lg���N�? �@�Љ�^���q=��:��8b4Q��?(��F�#k]M��n�N�rd��� �Y���:��.G�
_,ɇ�Q������)����Q7v�0c��¡�۹cT��k��*�'�l�j
|G���Յcw��@�A�J��L'|p�V5��H��7.=y�s����]�.�v��Ƥ�dk�'�#��C�����⃦x�8�oj�߅1�Aݺu�O���˖y�W��2�= )�ݶ�j�(i* �D����o}'�7CF���j�bg�