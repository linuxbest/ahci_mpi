XlxV64EB    31fe     de0�P,�'�%u!�	��_��/��Z9���팥�&_Ԋ��%�ʒ�G �tj(�fo��-I���*���gA�:NRotMܓ�ȡ���\���'�aN���=�ib���H����w��tN~�VOb�ᦸx�0�N�AC6a��ٰC��@P����e�퍲§ܺ��5n���f�Bc�L��"�6>�_7�0�{��佲�ZE�B.���6�p��iQ��'7���*o�(��Dg�WH������g
�����F`A$|�[�os�$�|tM)��ԩ|i t�_}���)	m��@�h�)i)���8�)�:6�E�����m������R�K��Q�#J��D��R�V�	�FZu�_$� ��u�w4�d�������f�񬐙��B�&��Bi���3V�d�2,y6n�/�dJ�a��I�@�z��k�~����f޵9�x��;�R����v)��+B�V��g���?V�HyR�7o2Y2	�����_v�%�3��'5���# ��㐮��4R���b�i)����Q���-4��5.��r��n��N�d�`�%�v!��qr,���R�e�4WU��@ǜ��y�>�@�+|l���(���s��ʽ�4
/�ַr�dYŤ*��6�+�j���,x��S5j�4�ҹ\M����Y���;@"���7'u��G���^���+�=�!W���DXQ@�n�K�D�p�A�����!���
�o��]/1�Z�T9jD�R��=v�_8����q��i��ѓ�l���d��&P%����2`:�`/�q���;N�{��Kc��?�b�/�h�%�U$ܜ��`�~:a�����Nα����m����F[޶��簪��Wo�9����20��W@�`�j]�313x{>y�a�'��5�#�MTz�+ |	�V��j^�DIW���|� M>C���[�2��榺�#{Wk���������΂U��j���2�q�s��r�_����p��(p��Y@ح|0�J�?;�#K����tθm��)�>̏Th��0����[q	�.H��<�;:?_�� ��S�&�O�Rӽ�u�7f0B�.Ww�D-���� ���$#������3x��K�$��?l�/��E�A�rƴoG��2q����,}sӯ�3�<�N� \��S���>�u,;��k������&��H��C%N��A�s�C&H���{:HO�	��V�5�P�N��^� �d�Z�S�y��a�O��tbz!�1��K����[}��E�,�j#c;�?1L�Y���O������s�J�;t2P9]���ap5'غU8B*3b���B}O��Ր��P�3G�&�`5�zLl�֋	�Z&�*��k�E�2=ʂ}�bJ-�Pߜ�r|�=��=�)zÞ���ۡ˪x��g#s'�m_�>��d-�E���z�I�zB�.q���S������N:"TͿS(r՟���ɟ:\T�vء��)\�1�n��d-�"���e/SR��n����B2���G�
u\A��C{\f��[��!�)DH���韴W�c�rj�,��pkR�E�&�3U<����@��O������O�t�3~��R��`��A|ͪ��ݪn���ˏ�F�L:��oU4s�Hˠx�+�ӣ�^S���H�q���x�i���]|���c�W���!����Ȑu�N���l������������5=��o���M��X���+���n>4)4*��y՚mp8�g�e�W�� a<�_an�MȮWn�`R:6j�Sö�T��d�����Ԓ���w1ƭMk�����ک������������Ao$�zl0Þ�2�����Ʋ��-uzH��H�NF�)_��	�a�p�.��ge�� �} �=t����S�f�7#	��a�깅��5��5;�7s?xP5�ZaLU+:���=vZ�J��/��-	��Fʽ�O.]��wYȳ�m.��L�.�_D�˪5����#�u/�;YK��aY�l��H���򩸍&+u�-Ai��a�BJ�,_�B@J�vV�]$�OMJ#t]2�q�nQFr~�k�-�Z�	�v�I�����G7�:�E��߅(˰lE�#���* �!�f��6G7y�:�P�';>�~f���(A�?�*I�!�����N�?���e=������Gu9 +��i���nX<��o�%���#U:�{�݄pEFhTb ��1��% /�~M��*�f�����juݺ-�֓���[Xb�۪i$�}�����mr��"L'�+�]|�auZC(\ r,:Ԩe+���	�aJ�5T
�J4�A��B�VT��4Mo�G�.�T�Q��_��-sB��T8�hş_V���C֨��W1M� \�k���*�Rg�^�����O��x���+���R�g�4+�U^��[����1��I؄����`�C޵়���7��]/R��o2�x��>���\��p+ӆ^���}#�	#n��*��<E>�g������f�L�� J��J�w����&��Ɠ�c�I�~�M>��3�L�\#��QW�����q�qq>�{I�^�
b�e�(�t18w�#�=�t�9�ʎn�ɮ7�`��)�����V�*[U��FZHW��5�j�ŋ7N`K����:���
��QD���	���ٟ�'�^k�R�N�������f�ȳ�J�����6�w���_�E9�4��8<�[,4ƒp hJI�i�|�u��z�����d��O��DQ�W�'��|ˮ�%I%`=n�F̛v7*�{.�(�R �%�KK
�����T�/ǡXse�-��n��i�/#�� 5?0D{���Ƃ��L�����D2-�Ś�s��`FY�"�W	�S-�����s=b��� ;�#Y�*P��ly���Z�����?B_�¼>���m���R|��n����>����)Cދ�,��Yѷ\�	�>.��%It9B⢡��R���d�>��[��G�L-9)����,OٌK�
)�^��j2��>�-�F���/�Y�M��;^�M�K4�c#J��pц��˶�Wʪ��rKbG"x��7��]-��k�x�fW:4���|��9̎��	t~#U�Nz&2nӼgF,�$�py��DR����_�g@	>?I��g��y��m���AѭD)<�Ʌa���v���:�ʛyW�7��I�I���nΖ���N����5���E��ؾ0b�,�\���	���y�Y�A@�T������O��W$F#	p��h�v��c|�~Z&0���b����mv_!TO�N�d��	\��4�#�~C�s	y?�ZB�ڤ-��o�Z�h��2�+���Y�^#��0C��f�����'.v\u��,�T�R���0�#5� `�n���  U6Ln;_x7fƩ�F���W��9�G~9*�*s����Hfqdr����8^�`�Yvr���w�5+����D��S/��`�����ɏ��@�^A-L#+*q���@��