XlxV64EB    8c69    1540���!�/���34�	G�V�3��>q�E��mH]�����uJO	�>MXK�ۛ�7�˔J.�Hf��P�uc�d����zh��@��Z��t6G/tmm�\mFu:c��d�H珜�ʎH+�*�a��v6h�N7�]�ڡ�-��gy�O�3���Z8�r��P��zr�c�%x�h�u�& "��ȝj�.�<r��i�|��0j�q7��^�˅�B�����3�:H���tX-֖n��b�@Pa���~�h{���I��&0Pw�� ,�)K�F�[E���^j�� ����� �#�4M:���I����1C�}hd�sj�Qً�\Е��I��S���u�+����_�ԿQ;�E]���\��ᅱ��U�ڪG<̶�Z��,����B����'5����d��3����j��������k�W5}���а�4m������_�h��E�և9�Cn�+U�`�
~�F�
�8~v��J3��>�{���/��j��l��#[)ws�W3�PA3SGR��c����3E�a���F4��R��ي�e�� �/���V�h���jqw�
v4��3%2Mz�N���b��Bu�W����3����E��6�3�|a0WJ��8m�����4����y�$��܈�H\_��$$��,o��w~���TBh0(�L��G��Z�)8Ԭ����Q.�r����8�����l��:1��D��Ձ�K+�G����D���	���J{�(4�cIT�2�߰��g�TPz�.�Q��A��@) �!�3�!��L� F3;�[" i�%m��gOj/b?!�J����l��f0�rL����7�38��} �%;!&�II=�|t��L'���?���˔����ͫ�R�c�C\�a}`1N0حg9�&x���	�Z)G�����o�7�W���*�^�bGǌjK�7Tw�~��O��z��� ��yc�7���f�<\��@%qK�z&IR��,�S�!g1���� O!��B����>�@�bF�[�lV*����͆};���<��������?~���5$0�����? 6��u6U=�M�W������ѡ|�1�qB��h��I;���5t)|��>!�!���^�Eg���H�2/�}z���}[/��J;=����F>�8�lNWV��i@¬L]'cyll�����u�@�4�`"�"�:���[�P6���x:a�&��Pɽ6"g�>:��Z�#�A���uk�4Qbb�!���ͤ�34�p{5�~M�/���c6��D������ޅ5L�$�"�j�ϐ3�(	g�ѻ�w���e�(�
�F�[���fp�g�p�b��q^����E���BH�*�1�� Eb Qɿm��Mf����#2���5��\��2c��6�	U�2\�����(ҋL�E�/d�B1���-�ʷ||�����u���]������ڡ!0b)88NLęL蠭J<+!v��ƅ���|s����3�؎�X ���$�Q�r0i�qr��?�5��b�(O�8�'�)Bfi�r�&6��Ƨ�>���w���ǡ�W����L����۔ψs����$\m�NXQۛ�7���nkPV�(���(O�c�W�o��	?�Tp��OIYxj� ��ָВ��z1O�Ց
'�^��%y���(���$i��[2���e��3����\�O���iM2厙姿��1�84*x��~�=�����x�Ӳ��
�GY���7�+i�[S���٧v,�=1���(�r�i�Y���_���ߨ��-��֘�)���,���s\�xqz2~�E����5Q�4�����?ϐ���X|u�)�m}�bm�n�k�1�W[z7�{ĝ�~摱��w"������J=����Hf,ǒI��~�+w���m���&�j�n��ҞX��"<��Iԓc��+���p�'7&��x&BB�}�q4MA�Ya�;3z;Q�G���Z,��
t�C�gWTT��//P0�wD���{H�Ta����)���xZ�vG��5�[�#z5�߄�|	1��;r��C�x�]��=����'��M�i����A�v�de<�Fi�Gj�^�,O�i�o��V"�E����!L{���#�����n;o���L0��E�H�� ����U�9Q��!�򬖘1=+��9}��q'�SiHy���X�|VT�!���!�GF�Gb���c�j��0_n�O���J0�f#.�
�2���(�ǭ���q��o����b�JT3��<S�>�o��d�4��%لe�/��]t�a��~X��Y3������e0��}�mѩ��9�yV�%m4����͑qu !S�i��9�(��z9cȬC��Κ��W������@�V4�8�\���L�FaF=uw�v[?9}-Z��h�����5d%j^�U�/�դL-�W\NI��pP����"���*�'|R�̡){P��Z��Yf���  OZ�nn�QǏ���K��p����*�����f #K�գ��)�,g.��p.p-���Ƿ3��h��1��S_�$���a�&	�i���I<D��+~�[��͙��2��`"�ӎA���ij���,�^�O���H5�#��6����"��L`���*z��d�t"<��l�_Ԧ��J�R���?;?]����D3Я�,4�ӄ�-�2�	ʿ����V�6�v� ��X!�i���ߕR ]y��ە!Ð�l2���2����g�����L%��'�|CY��s<��#�(�Z�z��Jv���+	���^��m�/L�y���;�{����O�Ю��$�5@�2���*(�L�4 ���~1`hw��̋*��w��^ ���H�z�͂�uL}f�"���hȭ�'jZ��(�����S��K�`�3I2>�G+�j����fCRf���*X�?�.�53�����{�l�y��{g�,�JN:��AI���p}iM_�o��qؠ+oV�T�bi*� \%��� �`!����Ɛ.Bh"�F��p?hyI3d�H�O�C��/4�$�*�T?���錗c�&o���z_�B����|p���k��q�}h<���k�,�]�
�<��44T��7"N�����2x�HmNѮ���M����($rE��mh�|1��q�0�WS�_P��55~������ݑ�����7b�Yo���d!��y�
a�1ⵍ�)�`�w�1��'�gǓ�����f��nϘ���)`o=�c@6#:8�S6���o�:_�Sw5��Jͨ��:��y�|��7�E������Q]�&����q�N � G��@��t;I^���#���/$�A[�6�����쨾����������N��)�)���"\�� ߖk}y��_b�2S�&!�f��$� *�MZ���FQ(���σ�H�#��	��@�5�5@i�s����U�W��GL(��<nNv�:��]��^?Uo��W;���� ��K!��:�ɘj%�G3�C?�4h��N��j�C����f���V �#���)�JY�ڂL����v��K8�H5Z;I�\~.d����9)G�dk�����m�@���^s��D׫�ۙ���i�,D��yft�-��%=~���xT:]��=mL���.����E<ߦ��Ԓ_77�x�5�(���fAqe�LR��Fl���h��pk^%�l���L���F�}R�u�}k��F�u�`���6�o����j��)�ѹ8��e;������ʵ���D���<�����b�Ĕ�h?��@a}3��2�*u�����w�-�.���G�NA�{N�����:�Dcz<M�6dL����Q���\��c�T�������6���7�\'	�{�,�}�N%�^rN�� �D�6S^nȦ�}I�E��	?:��;��ef>|9��W���i�߅>hp��T�_�۠?XSV2�a���@, ,�_�ow��y���F���
Zˀ@<�K���o�v\�/XO��]U�>>���Ԇ��9���2��X�(����YI�^F���,�8m�> ��pkb�	QW��4٩ҸS��sP'�3?R��, �XY�M�����t�NM�q.�R[S�%\�/m�k�S�vI���?8\�X��]�9�1��5L���{{��o}%��*2�Q��H�|��Q���["������ڐ� M�_O������&Z�ǽ,O��l%T���84tNPO�92�y�:\��D�������[zU��|:<�ŋ��e��>�V�)�|w�*��e"��
�x�S��a��|�7��*��8�P��P�'�,�ńR��Rj9�[s�Y�q�� ��-?G3�����wj���n�W��ck����l�IA����d�Be�%��5թ�9g�kS���a���{�j���\|rh�����ʉ*__�B��:�y���PU� �)'h�9�Yk��v���W٧�g]�[x7�k,���E�mf��
�~�qm!��JhO�!��>!IlΪ�t讶I�,D}MH�S�J��b�L(�Fe�nL��P����1�H๽����'\#��m2���P����5��µ��Ӕ�8�����_��'�dp���Ɏ@��4_�E�Y�|7:��+=�!��G��Suy���'���(����L7f���L����7-ցY'w��䆖>�H.�6M� se� �'o�:m�se�~ت�����~Y>��8��x�'���"�K�ao)}�9��[i�����J����>X�᳤��6'ޚܽ_�3V���R'6U��_������8������PCq�H�q�G�SV5XV��
!~�?C�@�N�b��5{{= ��x�Ա=�q�^2ژ	�qhH|�5�R��k2"��K2>��@V�-�z��ũvC������o����֞���C ��<��cj��T�sz�w-���ݹ�xPy�]����d�S�*����4�)��R�gyg@X�L�ƨ4>���<��\�<`�6�Jg��W����?�$Ȝ���"&Z^�� �mIL����P������ˁ(�u�YH�l�eV7
��qD;�[�Ë�6-A���i�w���ff.���1X,�|"`�7�l�׶���I�a[�V�����#Gvf��P��X�i;�C�_� N�γ��t(���|k&8%���s	�Fs���WI�_G�A��4 0�V4�����xf�4Ӧw���k=���a��.W����O��6���]I��g����x�u(����Q�_(o,����Kb\&����Ӕ4W{��w������p��ՠo�V�)�v2�~<���T��p�;D����F����z�/`{�1k2���g��idA�)ʇ��+ʨ-ȃ�P����`����_Țe�Z5j�_#��VN'�f}:��W�k�F�Jw���$X��i�ak��:WJ���	���$�&�������`�V�l��