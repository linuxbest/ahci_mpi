library ieee;
use ieee.std_logic_1164;

package lmb_bram_16k_loop is

-- BRAM 0 in address space [0x00000000:0x00003FFF], bit lane [7:0]
	constant lmb_bram_lmb_bram_ramb36_3_INIT_00  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_01  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_02  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_03  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_04  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_05  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_06  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_07  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_08  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_09  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_0A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_0B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_0C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_0D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_0E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_0F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_10  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_11  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_12  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_13  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_14  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_15  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_16  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_17  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_18  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_19  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_1A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_1B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_1C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_1D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_1E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_1F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_20  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_21  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_22  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_23  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_24  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_25  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_26  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_27  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_28  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_29  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_2A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_2B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_2C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_2D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_2E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_2F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_30  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_31  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_32  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_33  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_34  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_35  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_36  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_37  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_38  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_39  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_3A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_3B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_3C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_3D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_3E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_3F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_40  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_41  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_42  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_43  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_44  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_45  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_46  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_47  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_48  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_49  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_4A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_4B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_4C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_4D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_4E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_4F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_50  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_51  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_52  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_53  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_54  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_55  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_56  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_57  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_58  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_59  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_5A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_5B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_5C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_5D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_5E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_5F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_60  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_61  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_62  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_63  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_64  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_65  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_66  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_67  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_68  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_69  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_6A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_6B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_6C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_6D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_6E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_6F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_70  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_71  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_72  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_73  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_74  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_75  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_76  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_77  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_78  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_79  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_7A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_7B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_7C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_7D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_7E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_3_INIT_7F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";

-- BRAM 1 in address space [0x00000000:0x00003FFF], bit lane [15:8]
	constant lmb_bram_lmb_bram_ramb36_2_INIT_00  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_01  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_02  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_03  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_04  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_05  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_06  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_07  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_08  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_09  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_0A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_0B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_0C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_0D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_0E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_0F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_10  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_11  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_12  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_13  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_14  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_15  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_16  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_17  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_18  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_19  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_1A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_1B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_1C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_1D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_1E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_1F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_20  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_21  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_22  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_23  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_24  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_25  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_26  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_27  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_28  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_29  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_2A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_2B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_2C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_2D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_2E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_2F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_30  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_31  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_32  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_33  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_34  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_35  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_36  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_37  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_38  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_39  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_3A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_3B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_3C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_3D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_3E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_3F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_40  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_41  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_42  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_43  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_44  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_45  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_46  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_47  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_48  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_49  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_4A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_4B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_4C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_4D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_4E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_4F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_50  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_51  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_52  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_53  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_54  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_55  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_56  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_57  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_58  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_59  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_5A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_5B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_5C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_5D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_5E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_5F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_60  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_61  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_62  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_63  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_64  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_65  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_66  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_67  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_68  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_69  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_6A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_6B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_6C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_6D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_6E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_6F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_70  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_71  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_72  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_73  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_74  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_75  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_76  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_77  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_78  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_79  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_7A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_7B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_7C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_7D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_7E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_2_INIT_7F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";

-- BRAM 2 in address space [0x00000000:0x00003FFF], bit lane [23:16]
	constant lmb_bram_lmb_bram_ramb36_1_INIT_00  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_01  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_02  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_03  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_04  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_05  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_06  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_07  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_08  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_09  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_0A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_0B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_0C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_0D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_0E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_0F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_10  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_11  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_12  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_13  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_14  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_15  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_16  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_17  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_18  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_19  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_1A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_1B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_1C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_1D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_1E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_1F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_20  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_21  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_22  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_23  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_24  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_25  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_26  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_27  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_28  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_29  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_2A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_2B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_2C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_2D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_2E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_2F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_30  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_31  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_32  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_33  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_34  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_35  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_36  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_37  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_38  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_39  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_3A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_3B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_3C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_3D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_3E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_3F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_40  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_41  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_42  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_43  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_44  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_45  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_46  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_47  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_48  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_49  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_4A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_4B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_4C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_4D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_4E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_4F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_50  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_51  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_52  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_53  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_54  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_55  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_56  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_57  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_58  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_59  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_5A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_5B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_5C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_5D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_5E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_5F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_60  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_61  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_62  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_63  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_64  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_65  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_66  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_67  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_68  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_69  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_6A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_6B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_6C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_6D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_6E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_6F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_70  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_71  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_72  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_73  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_74  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_75  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_76  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_77  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_78  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_79  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_7A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_7B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_7C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_7D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_7E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_1_INIT_7F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";

-- BRAM 3 in address space [0x00000000:0x00003FFF], bit lane [31:24]
	constant lmb_bram_lmb_bram_ramb36_0_INIT_00  : bit_vector(0 to 255) := x"00000000000000000000000000000000000000000000000000000000000000B8";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_01  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_02  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_03  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_04  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_05  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_06  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_07  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_08  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_09  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_0A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_0B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_0C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_0D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_0E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_0F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_10  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_11  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_12  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_13  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_14  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_15  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_16  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_17  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_18  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_19  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_1A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_1B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_1C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_1D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_1E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_1F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_20  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_21  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_22  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_23  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_24  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_25  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_26  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_27  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_28  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_29  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_2A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_2B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_2C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_2D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_2E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_2F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_30  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_31  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_32  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_33  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_34  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_35  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_36  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_37  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_38  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_39  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_3A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_3B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_3C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_3D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_3E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_3F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_40  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_41  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_42  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_43  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_44  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_45  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_46  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_47  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_48  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_49  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_4A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_4B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_4C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_4D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_4E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_4F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_50  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_51  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_52  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_53  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_54  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_55  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_56  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_57  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_58  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_59  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_5A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_5B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_5C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_5D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_5E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_5F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_60  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_61  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_62  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_63  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_64  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_65  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_66  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_67  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_68  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_69  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_6A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_6B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_6C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_6D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_6E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_6F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_70  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_71  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_72  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_73  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_74  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_75  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_76  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_77  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_78  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_79  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_7A  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_7B  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_7C  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_7D  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_7E  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";
	constant lmb_bram_lmb_bram_ramb36_0_INIT_7F  : bit_vector(0 to 255) := x"0000000000000000000000000000000000000000000000000000000000000000";

end lmb_bram_16k_loop;
