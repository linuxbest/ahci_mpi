XlxV64EB    2444     be0&���%�Ċ7��qe�TY�s�TE"����wh�܏`�h���O�L*PNb�A� �%�Y:Q�~�0��gw��ļ߫v�)�V��j���T�,����Vl,�5z���O��iϊ�\w����8�2D�y��.rIP?tc�����+\3�⮢�8�=�;�"2c�H�)v�N��5#�H���CD~���oH5UG���:w��������6�.���	�!����zzGbp��L&���v�����Vl��q5��k�`��������ф�=}�3ny��Y�m�J�"�hK�f��욑���kq�G�ҟ@b"��6X��`$�)�����([���H�=`�i��B�}����(*���8���.$�> �܀m��|�n��R�;�$�u[��j�'�U����B�|g>��NB,�6DU�*V�0�S��\��� �����5�VʯPېCא�]��к�`=��uˎ;�	f��n�}����}�D�( B�iܘd��c(q�w�.�?
q�0�\�(����?��c�;�����>|����P��U�tT*��:N���f�D(^ ӡn�49�
��KC�G�=ӛ�Y����@��\�(�h2��m��/�L2P��U9|��B�#3f�a�,<�+a����'�����5�+~��|xdp�^�|�.���Z�ij������gv[�Nq��s|:*�����l�d��rռ���9?��c��'�]u��g
�3'��*̋F[�yά���DTYQ�x(��|<T����?;��'"#̽�5��Nف��6�*�b�`j�B�3(?�>�y��%(���������R�x�U��9�^�:Ψ��9%��R�)b,^1��e;yH+-i[%O��:�/�7_��5�(��a�w\L�8@����/�X���<0�f�����3�w0r{ ��b<�9X{���3�WR��V+Ѫ��ڽ������V��Y���;|ۂ¶i����?���I2/��3rfO^W��w�����<mY�i�6��U�ȅ���|:�o ��4	l�&<����dU/]�K��T"�{e��N��˺�;��Fxl��_"�b<YƆh�U+NNȧ�/�+<��(�X�lh�����;m.�j�Q��T���#i��g���v|0)����@�Ɔ�A���*ful�`J���\�Iͦ\$F����=E��0���@�?���C��]f'(yvVY�+R��sht���n�ے��y+���iXeH�o�[	�bLu��A0�zY�c촙�� �7��0���򓒝�����h�ʫ�)ժA�ιk]�q"�-9�ˇqثj9�e~BI���S��]s;�����a1���Y�r4w�ې�i'�/�__���^�B��g�ق$L�t���L^wj�(M�`��u�}�Gڰ�(~���$���w�(Z��'|��|:pg�{Ag��ɮ�%E��|�"Y��ٴmK7��S���S���r�$����FM�6��������=�]BNQ�m��:�H�L�|n�z&���cm���"��|Q��c�����Đ#i;�ۗdv�
���/��c~���&+���Mk���=~B%�M:4Q��$�q���l��HJ���w��@.�"�ZT����_X����]�c�2���;�.�:�/�ؓ��1��}'�)�w��:��;�
��q �8i8���9҇L�*|�������1O)��Y�o =7U�/�b�[S���^G��J�㵴�N&`#�5��C͛J���7d̤5~�*����a�BP���C&d�,bR�Zram��,d��oUV|���Z���~:�1.ĭE~_����!Tf��snj:����ǿ��ϣ���pb�p��ҏ�@6��"� �U�t����d��Z6�C��E
O ǣG���6�t>/D�gv��;CZ���u�e��?UdRH����}ׄ6.��F�<����(���J�;ֆ��+�d��h7vZ�HQ���,9��~D�Tm�ک����U�2]���U,��_f-Q}B�Dc�O���="�[�?$���"�����T��N����5�~�f����z`{&1{U�ߵO�_�	j�	^��F��O��O��������Ƃ�{0Jv#M��;Ï^�<���<C��ha��\��OP2C9�
u4v�7���U���I
Lٕ�S���
Qhbȑ7|�tw�J�����EMt�!o�Ǚ
����u8M���!�ǵͅ���_����+������u�ڦ�FZ��x�t2��!ݙԿ+FT�G��Z�F�ۡ[���6�lH��� �`sP�=U�	;ޯz�&*����7II^Z	Y�N���$���Qkw��+U�'�Qs6��PS�ԯi|fI�����
[�jL� ��r�,?�-��0sܠ��³��_�:?�2m��C���Ǜbխ���,�X��>'���É�e�?<� �|��x�wɵ@��a �����>a��w�@W!==D��ZrH'�����CƬ�8<}{sa���}���#�]��[�F�K��O�R�S�	��zH4����[�43��!Z7i��R��*� b�N�H$�;�4`X^�[�ߚ���(/sr�T��"g_���m�݀G�G�R�^%d�2�Œ�	p�#?��M�f����M��Dr���ew$�K#fTɸ�s'�3�7\������ޒ7�@���J�/��3�¿l�8�t<�I[C�˛�F@~��<�
vaK�O�xA����cra~���mEV\�rk=G�g�t��5�K��n�5h��Yf֍�O��$>�ܔ�U�r6Y|��-�d��賹d�����`7X{����Xlw���a��(�tT  �۪���_�%��ʹ]/���iB���ӄ����uf�u��� ������E� ���b��v��a�/�XȰ��V���Y�O�'�32�$U(���mq��1�[�sM���O(!�_W�%5��**gD�����7_��c��F�c��qs��fH��ظ|�Ds�����qvL!Ɨ�