XlxV64EB    9845    20d0saf9����	������$I�ʹ}7�.�(��q�����ӛon�`.�X�9'Ѥ�S4z#A
,�z�I Y���#� Fk�l��}��:��� l��o��N��f��z����#���:�&���]���[�r�y�ߎ����b�#k���Wi-���
���	]�����>ݑ��L̹/v�(3�կ ��p�=~�n5���>`�H��=a���՝Rl�i�J)]e��_*Ͼ�V������hz(������x�pe�I9�+׈F)�[ZE �9��M����
x@h7��s��
?�U$@���(�z����Or켐�6��5�)�̲��\/Ǫ4���n����
"$�aElJ�x�X��lt
���(�dt��;l�C�[֜ZgV@���ƥ�g;}��!f�����ǎXY�^�z`)�#Ģ�=�X��O����($Lw�s��\W����� �^�q��<Fg�0����^E�r��-/Nf�?-��ј�!;�v�){���_�u+�F*�nKFA��y��8ml�Y�騳���S���'y���1�C�=�-���È����7W��-�d����"��э{	��;.����V�E�i��x�y2��7�������&á�W���)�.eu1��c���"�&ߎ��3=rf0�j��뮘�8bQ������&�Zy�*Y�k��@����b~�^Wp|�r�Y�Pn\�&
	[�&sy�[u�j���u� Y~xәc���?8pj��|N�ĕ8`)���S��7��ơS
m3��g�>aIU���g��g�� �5<.mחK )�ݬ�QY��3��H����W���\8r�p�7��b,t�M�(y2�v(R'	�7��c4�[`���%���5��X�?�!�6�N6�vߗ�Yh�a��p����	hbX_��
ӄ|�P=�Hf�P�VEA�^���s��[:h.\�NL��fX�K�����)sz@�8��-�Е������٣c,�̢F�/+hN�R��衡+�z,	���"��#5�k\���̉#o�1C��}P?�#f��S{�I^�B���&�E�xƵ�egޢ�U�W���},Wzk�.dDaF�S��>����,�_79�Dտ~Z\x�7�<�2�q3]|	�y�GE+|�)�=D)��J�C���[�A��$���
�N���Y� �rlܒj�h-+TxW��;���"����e���8��ɝ|v�R��W�#!��z#}�%�=Ϙ�\-}J�0�\�<o�Ԓ��_���;�>p�F�\\=N��:@�O�^k�q��W����El�[����OI�nH~�qh\���m��I J�$ZR0��R-_�F:
H+OK�ܳ{]Й���O���t]���y:��^�p�G=	�߂�
���Їqp���k�s}������%��j2�F��$�_	p� ��ʹ����&��Z�\{�994_���=�40�L�����5��@�<�~����ǈӺ�t�OH�=#�WP����N��,�}���ߓv_�n�!+��q�U�=ݎN�˫���oib��k�cދ�w�I���c专|)���DUQ����<r�z $0��z���z?B�w�K��F�?+���x7`�Ǯ.M�[}���	WO{���+���b4q�=_)L�4׍�l ��!Mp���[%�赉.9.W�ҕ8�Wˢ@��Y"� �����I�mS�2�,=^�d^}ym�N�p��l+��z�j�kIB\��J��� �1nv���[��=ES�>���АNIhJA�j �Z����6��x�t ����ہ�Ƃ��|�׃�w�3F���G��H�ig��%��F����jH���.ͥPa�.��إ�jT�}���l����✻�����L���{�5����zH
�lp���w"�>�$�z7!<J���?7����-ԏ�����0�Y�@/���4�^{�l}�=�D�	Y�C�଱]�H����]-C�S�R֚$���h .E+ ��H�V�k�kv�b���v��6Q0�@ekw���T�m<�����Z)����X����ْ��Yn��\��h��mH+B՗ڐƎj��&���=!*�Ń`qLfwgU��
�������sa#�cyE@�b�;�Oh���A3��͡����u&�Y:�FWW��� ���V�bL �R�@#������TA��C�6���j�Cy������%��,,%����G2 K����<O.��������n[ �XXF��9ʆ��uT1�mU�"�tP72�����r�%s�\m@^���H�\���A��/LY�����`�Zn2���@y���P6��c�H\+�~�qkg�eQ�r��zT��?AO����!���3P?D�-�i����(z�xZX�����c�q.=���y2,�U�_��o�j�剟]��]R^�_��q�����T�ނ
}#g����%8\�f���朦�'����Pg�gs=4H�X��wߩ�j� �\g�K��,�ך�,�	t��L�١�ɣ�M#r�)s����Y����a��|L�ĩ���_��2�	WSiMy��C��0k���
��Bf�-s��vnu�.�.�V�
����Zzǉߢė�����J+�s�O�K�]|�)�T�d�>���B�ɜ>S<�E����|b�N"
J^�¤]26&�P��儡�)u�9X��izZ�e�(��{U��#S(�b��LT�?D�������G�J&�Q��K�O���f�QS��U�P����ǃ����V��"��#�a�	HC�p���Ӥ]*m�j��f���8�2��
��9qt����	_jUrbc��B��ī&��k�Yxe�fÎY��Z�XB먱�ʙ-�L:���V����=ڞ_f��Rf1>a�.	�u�G�9nّ�1��п��-ɲբ����\��Xݟ`?�<|e�%���W��4�� 'f�{R���V��)vI^4]4:�t�ٹ4���z|� %�.�>�m��5�y�(k#�Wtn��|[w�s��waᵒ?O�^?t�!9�8���"aa�z������Z�-�b�Bf7��Dt�%��Y�q%]�������`���yP1@f?���[q������_յ�ڇ��:�TT�]��IUc�{�x��0�xLdV���%������ ���ڒ���QG9��j�(�W�`�3����
Q��! �ڊ�e�z�Sx<ea!��̌-i��Ѧ^�`��M�q�V��m1�̐�3�C�׹��9k�V�:����| ˞B�h�F`�J���oNR;;�}ފ[T��_�j�Z�q�\B{��$ �ZL,�̶Bw�	�+�4(z#������N�z'oq�t�~���Q+��k�%W���?�oM�M~�K�:jNd3`�봜$���4=�'SL�b_�J��k3B��W��n�X6���N�_?�#���О�x��X��IҪ�d}ύ�����'�L�����$�d֟����݌ɥ\�ױ3ZآT�� ����i�K�|�����h3?���{�Q�	����=na�<����E��g�E�>���G+)vg��:(r�����mԪ~�{I��wP�E�89�dJ�B�
1�Xd�Z�y�Y�#�����@���6{�z��-3��x��f�����)Ɗ[�]�J0uFa��n&E�{(;`�#��>Ju�:Y�8�7�+�D;�r9����p��'�����#�����F����'������d��B�(����OZ��Hl��v�
.�=wO�P�]�}f_��q�k#��4�l!kG�$�pz��7;ϾH�7��b�e'�&���W�o#�X���k�!����?W2��mR�pfvx��9�x�I���A;ĳE�$��L�7�݇ѿV˂�-P�^t�+��pF����� ��8nG��iZ�Wb���U	���g�c�7me92%�Y�)�$l�~Aq<�h��2���MSzE>k�/(�e4f��wh���}��d�.8<��P��<{��}�҇*�3�V4~��V�����]d�Ҫ?�φ�����`}��	�/��8��,�	��ߤ1���Am�7	?y���+k~�����PEȄ&�˴GJ?�@��z���c�`i�H�q��p^4��fYB	�_�J7�{�����ƳL4|�φ�d����9vbP�F����R-�����j E?��8ly��.�Cfvw�=��u ���&��+��?�/�G!\��$l]��#Rߌ0���o0��R(ں7-Q�pd)o��,��N=��[���gw���!}��D~��aR�"��z/��Fp9mKN�_���{��y
 �1��ŸCܵ�9��$^&bu���$�������,�]�t��s�+�'V��a�]���[��t� ����)�w)v 3�dx|��8".�b1��1�3�v�3|�St�*R����{5���:账7W�(���(v�#^�V�����\A�˒�q��q��[�K4�}�Oa����'����,���dZ�/]9x�U��OGI1 p\E�A�cAg��t�������;�r�C�s�`���6�R
S�Z5߫��E��L�A�p����ߌ�J��^��y�6�� ;xݛzg�.�w���T�i���9B�Οx����W���`:�U�Տ�ϑ�Ð��	#����|C�����=����th�s7 ��/��4��B����F����A����%���wp@svm�vI=�!��0�<6�3��K�2��$��$��s�B�^P5�="<y`��ؕ��I����bos�`��]˺�~��5{L~5�7 5�J���#�msS���dk�>7�V�X6	t�R�~����.�i��U<��՗U%�N��\.ښ:�
�[%~������+��0�Z�s�]��(8	|O�/Svb�sBGh�߼�5[C�m�Y~�Q���S�4��'s���[�à�.�,�J�L|`��=��˿���Q�A���^�^�`i>#�8��F$�?��\�۶rk���6#6҃�;�2E��^�|y?R��?d`���.���8�{�+<��~ݻS:�Dעf��/љI��˟����8�7���+�-H��U�G����@�૵���\Gx~_D0n@�[��Xb���f�%b9�Ug(�J�~���Uq*�'KM�?����T�^�=v�Ň!���:���"�.��+��5� Z����ИJ
۾���Ɏ��S�v���d5Fq��RV�5b�&MoV?v�J��r-#D]=X���%��9�Gl�:ba΂�Ȁb)Y4�#���z�r����@8qآ�$�j�p.�D=�w��l�y��Cۊ5�ىQ�Q�XP�gxI�cM3���Z̓���'?6!�Hr��c�9�]au�iH�z�A���G��f���z�zL���-汹�
����<X�(�2XWt�4'�>;Kl����%z5H������0�F&2`��0�����(N���S�eh��$��1���bd�(�Up;��$B�&��j����TXL����t��Şe�v<�8&��z��XT2PU�<�;���(̶�"3��`�%�¦|T�۔w����\���E*�%��'���xx�B	�4�pa�F}O�O0���<`��)�4U�S�M�֦���s�0T>���}%�8&����F�:�:�����v��ʖ�SZ�������a�o���A4�%^��X��R3	��	 �px��c��~��5qSOח�~Aaܬ^Z�.�2�*7:!�`� "�;P"��z�)*8p�-��>����Ci�B0����9=��|#$]P����^ʎy��Z�P����S�g�b{@�֯��{b�A�0���`���p��Z��ǁ��@,T� ��CI�u�0�i�Hټy�C�~s*�m���݇փ���Q�}D�7U����������Co"��y� �4&Q0�6���H��*�#�~�r����u6�PU���[,�c�ƋEա�r�@	=*��Q�)�r�1;Ħ]���x��A����&ג>-���UA��}��cJ��3zhm ���,�z�m#L�!ϝ�ѝ�r�$��g�������>���Jm�G���ļz$c�b�g�vrq�-�G�;y2x�E�^��B���:�!��m�� S�*�j=,���0�1�K��SGe0B*1pW���`�"��l�7`�G�V��A���ڵi��H�tx*�h� y=�*�q��Cb��{�]�
�!X�A얖��3!K��,	ۉ-˒D^r-�E�l샹�S���cO5�'�GUq����I�n�����aI����y�k��_��luE�]?CU
�$�"����hJ�̈�4Z��r���`{8��h8T���b��*���z>��)>��2���5��������K��ǀ���S�CL�fm�s]ʚ�	MV���R�E�Ĉ���f�pq�&��Q��5&�kQ��6�����	jh\)ؘ�o��2�5g/�j=azF�|c�S-�����ᰢ�ć4 mR)��f@�Z�z�G0���r��@�3�p��M�0����0O�����.��u�JN ���^0ɇ6�i���u�?*��x�� wk��SP�^�f�S%0|�o���0�R�p�K����e/UO�X<���)t|��f����g��S��,�FѺǧo�X�j���ʑ�ͣ��	�X�V��2�l՗�+y��ބ�_eIeR��_�X�i_g�}��n.7�d�_�Q(b�h�`$����9�zP��6�<�$\'z'�ef�x���@B�A�G�X�Qb`�����n�摒ճ�;H��~J�9~�Ҕ���r[N����_T.QLP�����l���`/�$�q�ڽ@d�44������*V�����g�g��*�&���u��\�v?��y��W�k�����f�j��V7H��gsj���&N=��4m�p�;���+�dO�Z�ľ�3���³�dWܼ8��r3gA�C`����D]�[�-_3��"����n�{��û�0n���a���b���s���&׏~+�$q���}X�H׆ht?A�]X!�Ǥ�������?�[�ٚ�������1;�0�|{�?��H�N�{I��d��K�+�rʉ�َ�4hj��?�֭����M�E�{X7�g��~(�oEg:ѓ�t��.�4�L�)���i�c�њ \��!U�Ei3�
��{D�b�L�t��D���+�V�I�2��1�
��.�e�ːMۉu{��'��/~0�q�HI��=��PQ�6ˏDW}�n	�v�V��Jeݜf?b����!��&�^s���
A[(�,`щ�g�n���F���Ӏ���"�e
���8�DJz-��tP�cze�E���8��1)�\���>E��<�u��K��#J���?z ��#~���n���N�#�e|�Q�;t :���tFn�OY�k~�̓��Q�(��E��^,���W2IV=nz��n0�Q/�L �PV ���&�/������w�5 �s�Sb��r���U�7FE�g���f����Jң�C�j0��a.�i�y]�!O9i�H����ö�I0&�h˹�O&p��v�;F|�+GÍE�SZ9;�q�$k<�F�^3����4�d��Ug���4K��ߢ�d��~��&�]0� M����;4C�s�d��[
6�:s�x��u����z7��g�&�i��)X+��:�&���|�g�����譑��u��+��X**o`�B���[��n�m -��[krCm��#�;��s�[�0Q�adC�P�V&�&�0::+��%Ԗ+���gd(K0��s���&��p�:|W�����yǀ���Φ]X�P�[Ć0݊7l�Y3.�V�|�z����ut���RF��mv-'k��l6O<�>�"�x�[�j���:���g�?-e9c�� �`�.7X|��@��Jڔ��i�AC�~��i�Bԅ�m��azĂ	�J��.ͅ:WZj���.{��;�����^:�*��8����[���{����m���c�;I��i���N&�Bc��-Gs�,t�I=�?h�r��B,��-Q�0�XlV���C�a��s�����a@�*�xOs%P=q��F~��޶q��Dh�X��5���r����a�q����ϑMso��;'$Y���R��!2�V�Z�#�vz���,}[����Dy��흵��ھ�#��Q�'�je���I��;.j�=�=/�a �{�O��L� �wv���%�ی���X��^N�m���,��37��)Y�H}