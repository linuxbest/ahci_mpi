XlxV64EB    25b9     bc0\LT�U�V�M�@��s�ٟH`��_&��Ҝ5U�B��rd�U�M��&�X�H7(��Կrc=�� �H6��Jxi�}����?�coJ<�B�a�*R�v(��;$�����s�-U�q��pM񗽖����3�T�30��0Q>}���ŊE�_-D����.���(����B ��Ce��p.����ɳ�r��w�����Ƌ)������"�F�C�Ym�+1�E@:�!���un�.��6��[�����GP����x`���>\/0�����z��5Z0r5�:�ؚ��X]�W>��xO��
�7�ۥ��+�v��7jX4\!��4y8��QQ��^W�PnV�y��g�8�F�w$�=�u~[<�\m,Fɺo��b��#D޼�S{<�By?|�k�>Ix0�ɿze�50��0���Xo�p�7�#��æ�dU�ū�~�>쇸iR6�̉l���q���k���Gݻ��~�2���º�h��{�x���T)���h�q�V��枎�TiL���r$�D�w���*k�*����2ɪ�k�~�| �Oø�ta�k�4e,"�`G��R��C�Axl��� ���A�Ms|X�E��ż��_G!�V��p�Z7j�:�N���r��*�SyUqc�����B>�C4f�&2ԍ]�'Gw��2z���
6O���,u����S'_�-Z�*�5XS,�x���ҳ�h�m���E�ʋ�A�����]��9h�������?�zu'�|�d�4�fY��d!ӣ��^�_&u��>�L��9��@�mx|�Fޅ� �;�� v��^�>����p��Fmh�0F�]����Ra���	ۙ��PkY�B��&�5^�,�U��� ��:{C��`ZU*�����>:/�,J�~���JS�ې>���3����~xN�A�[%g���y�Ch��w���_���� @Z`��v�?x"S�,�y}�b[�a8\_K�v���B��i~R;w�Ze	��{Z�B�3�� ,d{W�b��O=yL�vJe���f[p�~K����1��A�Rkx{���C@��V��xUH���I��l�����oI���'n !�h�a� ^K� 2�IԤ�=YPJ0as�%�o��lQ�(�
��'̺���Ď����D���?���)�{m*QD@@����h�Oq��+d�$�TS�	��e� ��Z��2`F5Xm4�-e�R��r�Jx���(��8H�t�����m�Ͼ�;1��c��҃�ke��<�5e%B~@4��W�d�Sh�L$�v��D�=��U���3EL�]��*��*�a��V�kP���n����D٩�gw͒��aF��H��s_l7�&�p��E��].���S�T�D�(o!�9	oD `aY������:5��ϐ,b����$T���i���_^ާ`�� �a�T���"���dŶ��g�\{>N���/���+��҂��WG �ݚa`���Y���B^�b�Ap�\��_۶��Df�^�-eF��`��[5�.���(8��Wg�]�FG����3i�\���ڧT�R/@�E�YN���f����0���e��v�j�Ï�d�?4��[�'��dp"_��S��=�r�}7�\Zս'�k��Ft3�%�g�Ly�᾿%D�F(->�=������:��_+⌌筥�w`��^��k��,�O�AO�Z�p0�ѵ3z�#C��Y���Bn��iڟ�5�^��K7��uS'[X�1�R�Hۑ)�vT�� F؂ԙ{!3P�sGq;�%�
1No���L%�_4ϑ���7N��PO�z����b�/OETZ�N���c�ݨ/��,�X���4	Ս�)4ʪ��s��`��t��H�`Z]�:/��UA��T����5��w���`�M��E��߸����?���a ф.������Ęƃs���2��lDrD�Nt]�>/��<3VƝ��"�)��G��rxG�2� +�դ��������
�)x<;��ӎ34�E���I�XP�;jrH��sMS\���,��nK����k�S]Om���h@ީzq&�4������� �y��\J�4zc�#��h>��>��`�}������+u4��P�G��P���[h�������%�B�|;zY��1)�Ǆ�e)�Fĭ���Ȃq�������j���O5EΏ�D��{�HU%r�~a[�1�;��^o֎�^��g"��8�ּ�Ꜭ�4d��$�=d���u�1��
ٴZ`�A�-��vp��o_��1=�6+�n���gr)��T���@��-WV�ר��̋�X���>w$t�|�߂�8�����%0v��1��w1X�F����LgL��[��Q���/��x����%R,$�>��3�h���VX�o�s�Q�Wa��c֎�iɰ�\�?nC�%��W'9��)��KM�s���X�d�X��媸^�:mDm��\O�<����u;��L�r��%�ȁ���UMK��gfѝ���������BO�N�uc�oA|��b�;�d�a��Rx{�|�{��v�F{���R�g��}�?�xҐ��y�#��~y��(��~��0NnFQp���+��jv��-}-����p���+M�OA>�P>Q���������\$�Z��e8�hy��!r.���>Zݳ��ԧ7�(p�����f�/X� C~F��`��=�k�>��Ǽ痪J�6�@r'�;w�w�1�x�\�"nhG�k�q��[1�; �ն$r��Li�??�U�S��
����پ�FR\;xg����hg(�êmS8
���TU_��gy ����Dh��*�!5��y�hz�c!'q�L��ː[�n�9S|�M�+vhձ։�1@ݍ�
�U*�.A�s�~���HA��]�͊�W�ʐ�p�aR;�����G�+bチ���gY����n�A�?��mt�w"�Ya��U��w#K�����t�to�m+���]�%�X���T��rU6?BS���8G