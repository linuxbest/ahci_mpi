XlxV64EB    5ccd    1430�ݥ��.�Rʅ�T^��wx�����ό��YG8�yV*Gn蘔�t	֣�&��^����y�~H��x#�Y�2�o6����l�5E%�DE9m����Dգjj̿|��Q;�pE�/G��M`VM��A�s8ID'�� ��^�h;�����ǽd�g6;6��4K�B	�Fץ�^e^�%;��rǕ�p�O�{�P�R���:���сg���GJ��~� )���wW_�ѫ;���9+]���/�bJ=���]���كM��(v�ó)�����~Y��蕸uk�?`�/wRU4�v��q�z4<��x�s��)ԟ��{5}4wk���4: ��s�d1Oo�6qj��	d�w��Ex�O
x���5z���$R�I�8I:�*�;I�ڨ�M8%�A�,:���g�q���Qtd��v)�v�5>��j�����z�;���0Yq/���@�|�n��}�Oq���8ks4i꬏id� �4I���o�2��Jig���u�O*��~��<.Ň!��.�@M/V]�۠���!���ٛ��T�d��Q����{�܆fC�<Wq�"U��2�	�$��z�DFL�^�dha����:��
۳�U����MHDd���0H�(�m�P��>�c���zP"����]¨�^�'!�8X.�tԻ6�r�P�g�:EI�ۃ�y�I�R�23���Ty���B��ޟ�@JT�&��%F���eI<��Q��8ª)l��ENL[�,[���A)OV��E����Ql���G�e�}���X`q��ˏTvէ�H�k2}5�$b��#1r���D��މ�z{�����~S\��&����Qv59�
v�\42[ [d0k�O{��P`V�����7�P�_������K)ut�̵�b��(�s�l{T�|Uh���TP�`"d��#E�I_�t��
���qa�*F��xW��;������*����/�\4:0�V8/���YH	�&3���x}��g�o�ڢ���2�vN�m��� }}V�����L��t�O"�Iy/V.>�^��N��$��o���XpD���|�`�j���Lk�iv�v�}�e�>�zQR�hگ�O-�7Ë�hz�����ѲLѼ<Y�� ({��2	g��7�|�� ܦWػ7�;�Z���k �-�ҹ=���/��ўl]>���\�=C���; ��}P��3n��"�)����[�5�c� ��ݛ��շ�t�
A��r4 7*}����*��<Y�,AoN�0��\��6+A��H(�؞V���iy�T�ފKVy(xU� �L�!cotR6�ط�P����O]�o�C�L`�s�Q�qK�.a`2��l���jh����Q��^O��gO�t��p	��tIh��d��ԸJ�F�۞mW�E��gI���3Y|�-�)��X�GL�DX�S��������3��ګW�mb�#�/����*��%GX�*�<�-�|�������6�� ��W���t�!>7��[�qK�1@6O\�q$A���

��q�W��C|SZ~�����0)�j��lK�:{�Ʃ�`��+�j���U�GaK����	��+�i����6�k�SJ����v���*� ��p��UYY�S�m�^s��r[�󚑦����9��̵D�
���G�F��zEਟ"����wB��g3��R�A��=]_��I&��N3��㬈�]� �J��zS�J<��h;�Q#����(욵�����/I���G9�O��1n�%�)L�Q��ċ	R�\l7���e��F����dZ�V�|<L�v�S��1�Q�W=��{9' pI��*�o��J�>I];Il��2D�3rD�}5;���4��4�)e�N�����(��\��)��*6l�2��0T��\��< �q��~H�(� �F�꠽ڨ��0 a%D�i?���S;�c�FV���h�vc;k���9݄�m��bNZ�y���������q�p�&#^�0�O�H���`nư��A� ��K����y�}֝���c6#�6gl���q�S;>���햨	�}pW��h5^������6h�@�_6G˳�5U�I��m='��+���%v�X��bH��`an]�_H�A:�D���@c�n(ٗ$	_썰�VZpA�#6�IL�}5D�4��C2xd������r����у%q���Me֛�3f�0�N,�yX�*����߹��֘?�'Y�c0Ѽ��x"��d��>��@��j���&e �y8�.��k���T��n�+�9\���X�/��繌��,f�`�x���!����(x��9��
[��˃��P릧��t�J�������5������c����E���m�b��"��^38L��0�7���+M��b�����(�].���6TB�᎛	�Z���	�[wUU&|�#�m̈�$>�~s$tkąn����U���7 dT�!r̒�{�u)%i7
��P�	�Rč�Vٶ\8+Kh{4Ʋ<����� �\�������**�,��s��g�6Oo�SX� �C��
ĸ$�J�?��^��V�t��B6N�Gؔ�ު:���͒w1#���QQ�"��o����]V:7+��K���aBu���2�u�:zi�),�e@�uE=b���gz��H@ૅxQ�/�ͻ%�i�Pm��Gpd{H��T�Q*���|c����6L�`�z�ֽ��Ӿ�)'���AG�)N����H�e��h��)�+���M
��CͶT;mz@n�vw�o����C�G}�[U�l�����t��OrF��c�oE H�P�:?��d�e\b�u�dx���Ɉ!^L�^�N�8.��x)Vk�Y �5�'���BtL	:��l$�B�#8Gk�� 	�|8���B��X�����r�+Ja'w'{Z�U	ǀ�}}������z�̬�������8Eز��`�=���@i�<�s4�h��q�hй��&͛Qf�\���3%�vOH�H
��8��ɭօ���ȡc���xgk��o6���������"ƴ/�fUT���M%�V~O_[�����~/�\68x+9q]R�.��`�>9q�U���i��4��Eg�%�8͟g��R�^��^��SE�]��f�զ�6]�mV[�&�{�^e�����Ѳ���G�.7;��dz#��-)Ȥ��E���xjy��Tk��Y��3� �,��̬�a�7�G���֌˚�<$��W�v���_��x"�t���d�^ y�E�����#c}���@^A�H�5Z1\�ւQކ�A�����^y�}��+/��׆������<��)�Ɔ�"ӌf`�{F#\{S��ܢ��=�m�L��jJ�(�7�6�b�t��q���W�����q�bR"J��V+@L/��&�l廫h��*����&��\�mN��N
�[����!Q�WW�-e�
�	K��EcC �p���e�V�(�D1u�q���[��Kݗ��l��{�|�̗�>�E<-`�^����l4:I�x[�6����c�F![�&1�.�5}"J��ǚ';��[�����E�E9yB�N�U��0[�I��<=��g*�����e���p�H!}m�D�{)���9��R�(/ �J��/�ܓǰAnj-�t�̂
/h�E����Ȯv�'%E���1 '⡙x��ޞO<�"~'Az�=��u��T�c��
f�*̌��m%�͂�quw�D~ h�1&ݱF�ˀ����?ϰwem�΅R�Z�,��k�q�B�j�\���Ku�Ǐm5'�]���x,��JXd��*���/L��.h�\��/i���7�l�5���J�	Tz�/1pPlJ�ۤ�UN�.���S9�r[�x�б�m>c����E�(VԶC[�u.&y Ҷ��"��mŰ��[~xN�z��@�]�$�B3�Ʌ��=^��[-�Q$DeJ�X��1��_� �Y�u0Fg�
�
��í��e�X�zm� %�EG�-��5r�}�8{�)�d���"���Z2nޯ"�\Slcw��%�T�$��s$U���[������X����mյ.�I�]��5�;1'����� ��ū`A�o����>?��E��ԙ����|H�-�X�ӝ�AwZ�C�����q�]F�	���'+�93�|J�(>QAɼ���Ԕ�!��a��4d��S�HF�ɭ��Z2���L$V�~?~p=�d=J��Oւ�䃢ɛ1����������yټk,�>�:��3���l�Gĩm(��bt�|�(m �Fh�e>< ��C��a��6=���[�!싴(;���@mT�3����w�_���,8j�0�w5kE�=os"f��\�~��@�k�~�!�ì�+�T��e�F2�r�7�~M�Z�垿罖���^�k���*ȯW��n9�Y���e�)�t�roǯ}�dt������w��ظHm2��n@:UJ{߈4�6.�e5"�'W��.������T��y��ddӳ�������d���<p��r)��!L��Y�yCɶ=�q4������!��h$T��͞��Z6�G~�3��}ٰd��Rdŀp'�4����r)����؟�ƲyQ2��g�h	��|�����C��Q��}]����#��(��@�t��'��
��yN�5��(IO�G�t��);+vV�-� o���ۥ���We�3S�߈��;����4��\S	�\�T��7ʺ6���U���{�0���iOB�hY�m��Z��T�Ǎz�[�y*m����B�ʬ����bww0��1� ڢ����=b`$�ˉ��&!!*�=�E�0���M	f�z��s̏���R���ű�Z�S4=J�/��Hh�4��o<����F�Au*�'�Үәa3�&}�Ц�����W�u�h�>V�T+w�[A�ls=�DޔO��Q�ce��cJ{g�:��8D)N�~�C��{�kg�6���i�Įl/��P/�10��(6�v�[����9�-6��߳�R'���me�Q��S}H1�������� �ܴ�Jҧ�"�����u