XlxV64EB    c84e    2590��fu4G��
"��XtW2� ē�LP6�fAg-�G@Fh�$'x̀��+����9p=���nq�� �mr�fqZA�yy��.Zm�H�{�4<��w\Q�-ʞ��v���2�V���Ld�|���j�%���w:��ECL�rc3@�0r�Inx�RZ�6&.����}���	�MSg{���q�{T)6�)��d=��ƶ��#I�� %�Nb���MC�`~����&�j�4��] v�iQ�(i�_�Z�P�h|>��5�2���.4�g�2�h�H����co�еRK��5���z�i��S�V�?D�������Ч�h���4Ti�O�5K��<k1g���b�^�/��'b��5F���`݆К�a��bA{N��gr25FG�t~9�E �,G�u����T�G2?O��f���]go}�P2���ތ֟��������TxV��~�֐�7x=��?�ty�5O���Qz�Of�q��7u�;=��l��?g�5��kv9�w�PՓ�)!2l�&}ر��c��6U�F�K������L���⿺!��0����]a���,
���O�1( n�95i����Z�W穸�2|s���F��K��2�kǭ�v�t�fx�/�d�.��- U}��&aX* ������B��!�R�;�W����Pr�%oVݗ�p�}KBh���4[���\:p�F_@��wę��.��{"�0�U�d�aI2U���>�~�Ϻy d�>+�c(i������y��7u5KQ]P
��O]��=�0�e@�}wYkޭ�~u�GF�z-ӡ3g���Bcvn��%.�v��,7�1�*9��B,�l��l_���Emp[����_V�F�X�T��ǮM�c�
��@J�x7�b�LA� ���"q{%:c�N*p�3�l������HmQ��6�4�:GK!�/����fb�jȲ�vES�!q���.���`��OC, ��a�Iפ�S�3D����rPâ���Ʃ���-UD��"�#b�@\[I�ќԕ��l33ө�+��u���"��s}F�L��}):d�j�[�B)��(z8�}z�ڌ@˙���^�B.肒d�3��3�~��
�9b%�HA�j?���~�8s�_W�T���(�D��	�I�������Ӥ��1�K-l��O�"|6�ИE��!T�ZN�]��uX-*�e�vf�R����C��/��l��T�!�Z���@�> ��k�5Y=?�1Y3}�ث4� '��jx��R�T�	�¶����������@r�\ b�,��'�HkvSo�('��Jn�Ƃ�W����4���w�����}�!��uZ�p��	��t�w��gt<y�c#�a��@`;G���D!��P�0����p�H�3�=MC(d�����nuJ:��5N^zv�}�O�Cyۢ{S��@N��S�D5�ҫ��q&s��� ��?���Gw��ݢٗ�	T���>穂-Ae�������3�t����d�R��ɺ=�=��Ph �?�J䗡�[��;S=̐�	:�����
yPF�kH-�rek���u�3�����%0Z�s�1�d
 i�@�����iB���4z�g�>��u�[�7�����$�_G��p�r6�����h#8��0������N�|�M��$'3N6�Ժְ��e+��DKz�� S��=`�7�X�6���Q�
f�.�f#�����M�z^���*<�}ֱW@#s��hs���3���]�����ƌ=t9˿-E<��E:���,wJC��v� *E���p;=٤��Yw�|�Z�C�U�L��>X�� ����C2�\�7ƿj���~N�Q��9����󃯡	pp�)+uTC�T��0e�����<�c��#>�N���o���V��j�����I?�H��U�1vi��Q4%�D-���r	r� �E��#�����ȡ��~��wo�=6l&q1�A�RX��(	`��;V�B�:�/I*���sH8A�w�/�O웓��QYC��:B�F�Ɏ oʱ��Zs\k���ԍ�r.��Xs���Ŕ��D�r0,Q5Z�q���Jʌ�$o��򲢠������0%蕛��׎��J�[3�ͦb@H�8��=A���ǻ�l̽
��'��jŗ4�V_�(��Xuj�Xl��^wN�O;��I{qX;!�0.�](~��e8�����k��S&&�MTb��"	Rr��]d��]�ZF�r�^����Ue�o���b4�G�]/�~3�|������d�*W�(Q�1���C2��N@'|Ï�et���
����8���mV��Lr^d��=[��ʞ$J�z���[����������������h͸`���==����)�o�:�{O�/r7v{�n�ʫ��8����RT��;����I���jSǤe��"�p���o�h�������?�7�����=r�Db'ƍ=�������+�G:����M�ŔkU���o��+w�L��o��^粽���mP�U�
Ā�q�!U;oSB bz�=�xh��hb���d�.��/z�ѫĊz/�F ��P`t�ͅJ�9���o�'4��@�h!2]b�7/o)�S�)bk_s��o_t#	"Ei�w�ٵP�!�h�R!v�}��.��VV�J��ǧd�j�
��ɕ�x^q-�r�-c��F�!��o���CU���ȏ��E6
��'�4h�n���BL��%��Ty�7Q��������o=�/���,郆y+��xF���c��F�M2��O�������s�V�"P/@� ��íV�s��;�	y�m}��:���IL�e��$��K�0�D�t�abP̀4g
*!����b;W����*�d9q�v#��4�b�e�a�����7�|DJ��]��A!!fՀ�u��Z*����Lݷps�_[^�71�^����lעL{���Z�YYJu��e�Qm��aà���S���G+(v'��_p�L�nv8�U�.��މ��y��[lY�sÿ����e?	P���ǌ]4T؃3�qU��DEs�߼������ғLb~Ϻ�����f�ު���N:�:�y&��)�g�#��g��	T�F���z��
`
�bk�p�'�z��[�j�̮Vj�C�7�z��p���ҋ9G�.PJ����~�q�?��ˍ��'RN���b�B�t9a���w8F��y��l��h�_4qk�~��shw-��Нwl�.'X�t� ��K�-�KO��R�cq�X���R�8�>�h�6}l=u������J0DC�'� 7w��\�.�-f�I>6�8H'�\*��,/Ʀ9��9CҮa�?A�|ސ!���B璴4�72p'I&U\+�^5��К�ڞ��4m���N�����	�W-�<�zz�9�e�[xԷ'������±ޚ������_�2�{����c�$]x=��Ha��'�n���6�r���0���!TB4Utu��Qg���4��d�Jf��PA�t�,há�$�pQЎ Γh+<��|l�eI��_,5qT_jv�}��1�r����y>z�(Ο����뻅���aH�f�r�#�ֆ�r7�~D�m4ǠzO/2[����������vBJ��v^-}܀2LА1�q&�Ŧ�L�N�a�O�)���������x�SH��xk��*�wČ=eG
v�>F � m�U]���#��7����O��7�%�Jkl��V�!]�z�Q�Z5W�~~qw�I�� �\~ւj[��\N�Ƌ7\&�D+[EVM��U�L�X�K�?�t�j!4�pύ	u�,��I.~�Û)H�1o��i���b�ϲ��A��hU&n��r'#�{�2�d��Ϊ�7�:*��#M�������k�d�`��aIU��u��~�'��͝o���?�Vs���1�a�XI���߱�5�r����o��-Mg����u>
C�e��a���W�Qܝi��{z�5���n�y��޸����i���ӥ��^X�9�Ӥ��G����Fv�����L�c_����陥mg��C�sfބr̊��6J����J����uZ���Չ��mZ�@NJNd�L���pö���B�;'\=��ǜ-9��ԉ8���:g���7���K�������e6燃x�����!���%�DLIb�E�K�9��	f�!�C����}�7;�v�K��kGJ�oE��J�u�B�1�4���K78�]�I�����M{��6tD��f���|r�3��_Q[=&A���E�m�k����%=��g�<0�SLzU#"
:U[�k�:�=ݭ/�i]pj�$��זd�� � 5/���@�Æ}�����M����Bo'��։�� H�m��GW5���	�l�b�Ʈr�ns������t��	���98HU:��A�LּO�u3͗#�$��[��$��%�Q�£���E�Mu�?���%.\/֖b���Q�%���B	���dU�-��u�5����pL�i�a�Q���?vot+A�A�, Yr�~�"�~��xn:Pv㵆O�I!OS�\<�P2�}��l���R=@��o^P����¯�unJR�u�=�� �/P�8zB2�b���O�����ʫ�3���'�i=:Rߘ�0J)�D��(�A�0����������Zz�-�&�zM��W�Qe-�Ct���e�b�&6�Z㠁�o���a<-'�0��%0^���]c���T�ow�s�Ɍ��c���!�-�Jj��2Teg8��L�>9�9�+�y ��,Қό�#ׂ�k��Z|(�T��η����[v�]��4?R���㪬�ؼ��A����  ��W>�K��O������]�8���j��{�f��9��^��\TD&o&��"���Wٶ�C; ��_?
���33h����;ɇ���> �hE��E��H�d}�a�W�q'����T2�_�����?��V�`h�/�ǥ.,��r��*�hZ�+����ьO$͜�&ޜ��FD&����X����7�?r��c��2�j'�8��H���k4��C����~2�y��m�5T�<��5<�fm�Xo����x���Qy`��/�Ѯ�������	"�p��L��H���tHa�q��$�&'1�K�E����B����;��t�1r���t���H�֯3(d�A_T球I�+yw�mc#�C���Q�����'g*$LF��[\�z�"��]\�.�z��T$a٣E`���q�N�4��Q��g�y�4��b �%<���}Q�'�6OX�p��3��my��qG��M�|�X=�3)�ܪ1ɠ7���,D����n߇�G�\g�eC���cR���<K�R��ox�/�o%�V��vy�3�P��z�^�XΖ�?	h ���r�� �-uA�U�5n��1���^��*�����|0R~��%�J�`�z��.��D�\��t�YS�%7ғ����D�O�ے-v�0�M�e���זXγ��+C�5/���"��%y��(�1N��)�?3ќ�w\�����v.�9�]AJ�3u,~V�(�8��������H~��9��~fKam�����:�~��`*|�<i�{B��l���o�9lYz8"��-�
�*f5^.��V����UP8�����?Dk��.�#�Y䚳
o'	�}3 e �3XF��hmո��M{nZ�)��/ȍfl'2��0T�"j}t0/�1P\��a��<��	��u�B|�:m`��C�E5a�];�C�y4�6u��ȂXQ��t������gO�Ǩ��DҋI��Ȓ��8�Tz���aIL����o�h�W���H3��lÆ)Ub2�}����U�v_�ߔ�V,6�߉���v���§&��ܬW����օ}9�#K� �x���dL�K�:4L;�IΕ*o�����w_���D��_�(Hh�J�a1B�l����y�'k��{�(��/xU[g�J��2���lB��d���K��Sy�u��wޠ��D�����^8�;� {���,YQog#1)��*(�2W�^1.��d���0�EuJ���	��� �������T&^V��	����{5�[b���^�3t�\������<��nL*���U��#YJLSW���'��L��7*OÜ�R3�_W�EcI�cK♰�n��@}��=�;*.n2G.�I�fJWØ+%~�wfC��\� ��e�GmPIy�@���z�l�Iu����IRL��u�����t )a���W��a���^��G���cX�?_9����$�����*�]�������U)M��r4o,!OIƪ\?GhBC��K����$UP�
_nȣ�D1��`�����{-��;�x������P̥��V%�&rZ��$���K eI\~�a����`۰��)�v/7������;/�ʋ��TB-�=�Ô���4_��2���cm���9�]�ŀp��/��Ufi�"��Ĺt.�z��Ɛ�k�چ��Ia�K0ϋ h�3,�{g�+Z_���!��~������U�G��@5{5��kwcy)w'��C��`6F��ס�Z��\~aꈍ�O�y=^�W�� ���	���̀�*0��\�J���_�#���ߩ�.Z�J>ah��),�g^qIh��+�mm�l�c����I��7����ޜ=��x}�/ �u�z8�+�%{LZ�{����b�q�j$#G�؉��s\����@|V�iɀ^�y�x��K����r��n�xX%U�*�_۞��au0�������G��u��ia��2x�ƶ+�RD$NЈr���v�
���姠�����mҶ��+(Љ��anN�x�#F���,�M�"ݰ
<:b�1mW��PX�tEJB��`9'ፌ��?M'�@��Lx�S�f3���/�����>B���Pº�l��L�x��l���S#�.�����;+G>��֊�\��>�S�@w\an�6��:�c?5s�VG(���x���}�f�8�U��眽/��,����Y���d_���ݣZW��C����B�Ҧ�B�'���ώ}j�QIP�D�4����:ZoXj�8K+��+�/�o�����<?*/4v�������U�*_1av�Y�Y���q������sV��������+@Ht�M��;O=l�%�Mo��8ʊ�/J��󶂫�p�i���(%�s�i�ބ<*M|Kf��Ǝe_�Do�g�KXN���uG�u)i�R{��P�0$����!$��Y����$��j)�`���dͭd*�ׯ�x�M� ۴9S��Z:xp�����z�L��Ε�����摗+)M�!(W@(l�Q�|���X���G�%H���?��}�NPva�z@�)0߸_��w~���Φ[�oˉX*n�;c[��*Eq��UB,Ƣ�tH2�C�2d�=.�,�L/��eŤ'�&�72�� �d$ulO~��S�a0',�^�3��k�N;�
�~x�jx�t��u�.{���q[ks��4pF�g���'�)w��B(��'��h�!H���(��	y���z)��c��Mہ�ߣ�:r��q� ���$J<��E�:W��R끘�����1�_�B��P�l�����ѯ�R���_�ڲ>F�� Y�����p��Rq�m����xC����~����(/~��,�T�o�7Nқ�{�0�\�PRN�%�40�<����\�k��8�������� ��re�L���� k���v�Ka��ԿwY+w����!���$I()m*b2q�x�V����~��|�e��T����GV�F�><�-�z���Fv�;�ϴ��'�=��c�v�%�`q1��ہnٛ��1�&���H�
mwZu�n��K@�'.��oR��))�[LͯS�5��t^��c���S��A�ʃ�eHΥ:ߨjx�c��L�N��7M���<QW��^
�b@[�
n*��Gn
XC���p}�gg����`d�ʩ����d�q>vF�������h=�R�ڌN��o�����CG������OƲ�� uq7��a��s-ԛ�(�QQٱ\(g�����OF�/�d��,cÎ���/_{����c��F�YO 3��^(�	,-)o/����Y*d'V�^��%�����5�'X��Ҽ��Ľ�h�ҧn�|A��B���lK����ғ��S�m���~�_4S�MBnL֜���~�QO���8��i�
�Ԓ<�����TLRV�葈E61��b�������ޣ�:Fɑ{�iG{r�v��A�S����S}j�i�����[]�0�G���k�~�������Z��������L��+GK���yēB��-�5�����:��X�.V�Z���(����G����� ����yqM���W���_b��u:�d��Iő?Ðo�i�&������b�3E�?L!w�-�|`;�6�颪P�z��0P��̫�0a�,V	�߭PÓ|���� a&�I��jP�"�|�9	n��S��U2�n�ԃJȅd����ahU��������(����"2�-�ZYGP�_���L�'9�*��>��s	}����$���G_����p�4��$��wi���\���T��5&��{���ǖ5z����<r?�c~��b���>�F�>ڐUng���w���z�-��F~8ޗS��3��@*�O[~,r;��o���=�uE̳U[ח;Q�#$��~�~4��<�d�t��X7�T���{�����q������`X��~�1�L�#y?�q% $@����PM� �xV*���u���F�9P���j�.})p;�u��s�nX��%ן�u�E_'F<ׅ}�����p-�J\S7���O7��Id��p/�#$:����O;�5�����}�s�+s3�y��#K� ����hU�@ji������|�� >��6+7�#&6��;�9}d�Q��[��9���FFHfaϳ��6�i�Uٳěx��ؒ��SD��bA��;Q`nb�j�?N8/��C���Z�� �F+-,qOM���V�*������%Mg����*2�6��h]ʃ"F���Ac_=~�laD���A~D������f�؀�g��f����xJ����mߋ�=h�=�॓�k�S�RS��1Ƶ�D5�J���K4C�x��+ʍ�)�Ib`�p�?����^���⯫n=@1�c:����sa����7� ��&�i4��C����Ae	�v�oz�#��\��8�������<`�}����\����2 ��G,�[��U^�H@�����/��3��u��Cv�O�g����sC�Va��J�H��1�wH������n��s�N Kv^\3��a�at7�R��3@Cu!����Vk��̴vJ�������J�$�댋�բ�5�o�`e���m_"�T��K�~Ln�z�vY^�%QK��u�����!��m#�a�EXn) ��Y�mwe#�]���)v�>?�|M	�)ą?�<�]������������AL���ո`.ˤ�Ң:�RD�Db����fS�o���O�Gf�b&z�8~