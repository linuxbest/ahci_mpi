XlxV64EB    2b5a     c40<ĘJ~�3��=�D��Ԯ���������=���:����4�k�Z���Ɯ_�`᪼��F�6ģ7�?4��Z�g�Q�I3����d&խpn
�5��(���:qHwT5�vV��i�N^ *���a~4=lQ�"m��8g�*3%��xԢ���o��ks�?�J5�s [�u_���`N���YZ�\J���({$�\�z����b�=�*��������U�v�<��^�$Q����A~þR��]�bdpZ��ҵ_���"7�5��-���-*?��ֺ��Z	`ϫ�@-��G	_�犱�J,����z�*��9�8ĉ�2�h=V�C�wʟGO�O�jf�ހ
r���="������?e�+�/��g�"qX�|5����������<	�o'���酵��2�����I�d��Zc��Gߤ�+��-�HkA������ꁿj�F����m���r��;��Q�VFr��;W�ӎ8Y�*^�4d')�M���>s޳��ϊM�h�#��H�0R��5��!-%��0֚����M>�"*�Ҋ�7�N����G(7Z���#g�+Ȕ�{�"<!�N�va�����e]:S
���"�K	.\�4]3ގxݝ�嗼=�s?��:��x4��4�6�����7�)��IE��"��7��������ֳO�*��Snk��0����QcM��7n�t�5`���&���1PŨW�:M"xp$����G��@��*C��H/�G��AϵD|E��R�q!3t݀ā�K��Io��Kʱ�r%�ch:D9tԟ-O3\�W�NPa��S´XQ6OE���o�&�8����I����>�RI�K1��Z��n!c/�� ���-��̣�,O?�Hm[ʌ`�Ҳ��w�S�	0U�h�s#��Ȓ�z�)M�����9"��~Ŵ�:�)P`�mx+,�����.���Ob@M��;�NGٞ�L�T��_C7ϸ�ӜAX��Dj��m�[r�k8$��A����m��4�hCC̲8��FG�ԯn�7����hR���F�/�]Wn�y3"�k�����!��F��1��Sn�:�L�An��ɤ6:�^?�WƧҲ��d(�h��v9n��rKd8�!\V��|	!2�ȫl�a3=�qb�H�|B��g]h�A����#�&X齡}+�F�H���O��@�
���"k*�� �I���>��ƲX�$_���X"{�1��9�)�Y�	UE@a��7�ז���6#�Ғ6*_=�|�;�=W��AO�����5k��Xo�RGq2��g0��昬K��_�{��U�:ާQΘ����bZ�~5raz��2셌�D�Cx����K���A��F�V��Qc�-�Q��:DE�A`q,��O*�R�*y����9R�6_��?���DtY�5�/���q�p
�P	�Z�JT�⯩���odw>��l���W^�FС2�[��V��'ժ�Cj'o�RJ71#|DrT�q�Qr2�(�sORɭt��\urQwo���3�K��Be�Q2ޢ������������?쪾�g9B#�1�0���;�o`]n�I|9F�z=|Y=��Wo&���d`f�I����d2�gd}�]O��B:��i���6��\�$0���氋+��0O���TVR�ly�e�F!� ^�P�K�Y���7��#��Wr��~���e��O�l`�4�{xf1t�*C]y��_@)�Sh{ꐳ9l^˚e'��s��̀�t�M�6q[��D������孛�jA�/; Ʈ]���*;��S�gѧO�8��T���yZ�N�.�_��٤�-��Q��e?R�S��q���J�TrW� 	2��l����F����Ka:���W�U<���J������W�Zc�Q�r=�dS�ª����|TS�0��������03��+�w���t�?�4�&G�"j�O�TBF�����Ĵ]�៕-��גE�bx;�qq!�qJ�w}��H:�/s��w�N������u�P�
O��r�&o?-t �Ǘ���j��:W�Rn��m
�Q�j}�5<�H�S�G�׼O|� Ie�ǿ��^hc�sK3#������,���ā�4P�c�FQuJa�*ìx��`�������m���=a��a��B����f���2,�.Y7�cь����)2���7��2sO%�SǱ���_���
Y��>���L:���:�u
� L�nܐ�c<�to�͞�A�zϟF�F��4�4��x/��;�`��WEf9�^��w�;�c G.]�껊�2�K�Fq�{�ObZ;MotWCYyGV�?�U���Y`%ՠ�x��;��!��9���OHF����¢6�c+���H��7�12F��je���t�Z�Wdls>{�;?Z'�p�1���T)_=�Gv�-�Pn<������ȯ; �� FA�hZĪ́Wp��V���#�����>kL;-O�8�:�k�#.��7�3�S�k�BYڂe�b���-jL>�v%1Z�H���9=UZ���PwU��9B�c����gz��A�L6����Af4�FE1NHIn<ԋڣ͇��k��j����+�R@KŹ��찋�F�M��Ǡو�"��:#��ƛƓ-+x�)��� `�@`�t}Ϝ-���_e};(��nH��B�� 䜳��"�ʷ�kn�*m>�QMgQ�L�[U&�'8,{��;��~n��T���=˵Ϫ�Y>GILnj�;��n0v6���e����a��6̮����K��HF�,�m����xr���R�n��@���k=��pV�C��Ȉ���.��S�BwM%c�Bc�LE���8y+uK�@�IF��@�[a�1�aTX�e���l����C
�e��>��ayS��.YqUp�*������ȘOȦY��bjڐ��\�G�tO�ʵxckU����,���;��!(k:ᦂŀp�3��۟�F�7�=����Ir���;�G_�{�_�2���W��dK��l�-y��2i��T2Rs�A�#�	���6>��Iz�$(�dpP�ON�K�}�<Q����7,�&Uy}&���967PZ$ ��c�!S�c���KB؇���P