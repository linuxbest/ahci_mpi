XlxV64EB    1643     880�Ѭ�����f�W�<�㸸l�:�����RR���{��^u�&ة�R�M#UJ1��Q��YX���&:M<�	_XlKi���Ͷ!�YOGU�If�w����9���噑%s-"O*��(ԛ!�
��N�<�/���}�D��pi��M݇�KH��1��>ݕ��e�1��k�ψF��m�Q��w�^�^c�9D��H��?
��/�*̱���
Rв��3D�%n�3*Av�h_e� � ��'�aĪ���J��?u�FDBL��>Y_kIw��N�j�uF�-�[5�w�x��(���8��T�u��H� �l��Ԍ/��Z�vi���/�Ve���F���3�0�ɴ{�W�K��@��(��TJ=�a�E_��Lnd(�>��\�k8��(����v�ü ��^�4��7pՙo'g <=.w�	���������c{�ȥB��V�x�|�1�h	��$�[�0�pUM����%�8N�����3|z��Z�\V6zJ	�w���s=��9��{>�`[PbO5.2��^���M���+q4-��c�I�VUU`�>���0"<���96 �v�8�,h&|v���f�>~)2�D�WU'���!�����.��������aEuփN�G4��)FX� 8�=�i<��a�w�����~��Z	`��^"��xPD��-�	�� AD;�s�#|T� |o�&oU�C�w��˳IWW�G��#:���V:�c'��o�#�>�3=؟��Ֆh��I>G����3*��}����WU��#��p����,z��J�����@=�AsU�Cp��/���RF�G�3Y�륐˛��f,D5�/�'�Pel�`�GA +!��#�a���|L����%0��^�s����ѕԾ�I.V��4����P�W�#c�A��94���j�j��_N&�c�2|�bd�֯����|a
z��4��e�XF`�|�����r�<�3��� �;�O���Xq���\G�O>)�:���)�Moa� _]�
|ٸh9{��>��d�s�,<��*$))��v�*�ql&¥B�Y�)���(A7'4uw����T����l{cS��tϮ�c�X��q��o��1J�D>Mil$]3g<[>�j��_U�����X{P�(l,_��C�ad�(���ESsM#s�Ư�?6n^Z��I��ΐ��n-5kO�yV��7E*�F��3B,:�Zk��z"���K��2\6�H̤�|p9 �r�}P@�o��:Z��0�����ֻ�@�\�s��	<�/YZ�6�|
#op�����v�Op��rʙ��|/�v����{�#	��d*×�v~�(%�SJ+�e��:U�Ȳ�V��U֖ոMjo��)����r&��Y5T>!ӿ93�H�^��2UX[Fnu�er�����*Vt�1�6�9ޫ:�@b��l�ʕX�18:-�?Ě�����Y�S��"��:+�R�k����
�������,*��t��e�G ���?Q�j(G�W XR<���U:��K k�Y®8%	Qu(xfJs7SA����Fc��M�F8Сi2��slp~����G���!ΐ��'v4�HR��_��!�K�	���ޟ.�J��:5X�J6�f?���ᵸ"�;��X!���LU�T(�zl��K���H��d[2r�Մ��]��9t�_�*�~��m(��S�O��D�Юc��x��
&g���?��\pk+:�(��tOs~S��ı�'�mu O�[����eX+����(��3�n���i�UQYy}�EA6�<��	lh��u�u��WS	�W�h�'�c���fa$e�۟���E]B�["�C�=z�F�9���B�������m��L0�"�$�k�����OyE,�B��g:�1��|��z�N%�q��y��w,����N��o}jnE�<��O���8���1K]�f�/����i1��P��+l�6��H�;� ��8��z�a�n^��F�gyH�ʍvG�pGY�C}P���K�CT��5P^��l_��VW�j���s���0ř	(3`>��G����mz7.��<|v��'�L3`!� ��x�����0
O�1�����������ج<w�7� *��m?�uS si�p
2��@�|*�^�G��P�H�����p