XlxV64EB    227e     b10��1�׶�3̇��s���~����7�)؀�6[Q�{K�2ךu��r��W�5�D�'�10���[jo^t�2�1"�t���|��|���#�����&;��l
 0��H0r�q�}�ZyI�4�Q��?�n+��H�F�G� Y�|w!����Kd'~M�P�ȿX����_�m�VI@�{�9�M؃�^��y�+!�kg�g;*�-uI�l?Ui��%6=T��������T�=W�(�9d��꭭�{Q��q���:�s�fjd>�Xm��ZH���Ƙ�;�/������	��SCN	���qn��,*9q.��Z����/�щDbW�� 5�*l�]fE��{�@���u������<�E{��g�V�#�qNo�ɰ��[o>���S(-�`6�0k�pQNʸ��̖)pTdȈskN�OjsI4IANdp�N<{�qa�Rs���.��k6�T��:m#5a��a'�'�<-`�Xf����ž�,��6�!C�5X?h�	?��F����Cg����8���Biz�����*׷ެQCx�9�K3h�
v�e��	�s��j���M�ɫ�z��jړf���}f*�A~����fC���y�%���`�ı��;��׿ɽ6Rtˉ�;� = �z'qj5��_�H4V<�|pIW��bü1�����!y�L��ԩ锬�k�nU��Ά�eՀ��c����Kn[�O[H�{�C�x���s+q:1|o{*�L�j`���.vZ�RqJ]>�fM��E�70$!inI��������B�(g����G�!U@wJ�{���rOCq�v���5w�}ru��DJr�6К�Ӵ����0�����E�j�*��2�8�\�vj��ig��t�Q�M�SD�ԔT�p�(�0��oG)H��c�J�m���
׃I�'�`��7�'�y�\"��B�Z�ޚ҈q�.81t����a�_%+�����l����<?v�D¾b#B�J�;a��.N:;�H�%4ǩ{*|�C�=f�X���{>[�M�)$;4�U�>�Ҍ8 L����:�祈<u��!55��&f.�oL�ax��67QWP�x
:�SK�M��<�!65�fi��O�x���R	5������w�z����&}T��AE����M�"-x������Iү�u�I�)���X�V�@�; �]�4I�H������!�Y-�Z$�ʈ�h�.�-�w����?��qx[
��B�,�ͪ�x$�i+&�Ӣ1�E��������j�+��M
�힇Kd	\A�QEfт��r-8�������� ���� ��b#��0{�nɱ�Um�5�΄k�0c������
���P�Q7�.~fI���Ki��PVzl�{Ѣ��agp^i�'E�I�<%um��������vB��t���?�l��C<R�s��lm?I��3G����꼲B��i����'VrO;��)�A���3Q��MU��7�CP�lc��a�&[$�l��ƌ��$%��k��S6������3�d2@lDm�'�ȍ�YR�؈Ȝ�G
�1Y��M�y��\�*���#ZƇ�k�x%�x�㉽F�5j`[���Ē=�h�gD=7Q����eOq	�m���Ž��զ@���- �4};��)$�2�m�U��_����f��Hv����M�T z�:��<�@+��
�����5���[ꇋ�"%q��?�������(i��%�bl{ae�b[#���PX}$�=�L�=�oE,򎐶���0��?V�1�? ��v��}��wu؊���X�6#ZXE�q/>!�e��'��{w�
_�O��L՞�y��j��]}������
��C��>����o�/Dm_���L����zn���ِ�}�Ō���ә,8Gy�W�)�O�|�!����mtW�]rܵ@��?��9b�UAG�	6�#R�"N2�=��ڛ��p_.��OU�}���2У�J�/�/�Bp��>�3XA�yp�E�ۘq�Q6 �&���r�a6 ـ�B�*�*�Y�O��i}h2]<��~9PPƟ�V�����T��ܚ��������l=}JQV��g��E�բ��+�.�@l���0���� ��3�|�2���z�(+R~��	��펳,�f֣�4��Ϸ�7l2�i��e�n�����y�6r?�1��;�pmt����� K ��KB7L� �w�I��=\=��N��6��0��l� ��R��D��P�"�Ӗ��w�{(Q���)��Ӱ����F^$��!��u/�D�j抰]o��2����=���܇D}M����&M���zXG�e��&�:&ޛp�e���*[Q9m����� ��8���B�x�+�SL�U牃�ms���D���4�"�� ���{���D��!���'M=����=f
 07@���t������ʜ�CU����1����P�*<�'�L�����J7�w�ڠ���%(����s��.s\�(�
�[0�f�l�,LhjOe��o]
�*�Z���N �:֞z�����b�3A<SD���Wɛ��f $l���Fs�cK!��T��+O�S�ݜ����h5g����G�6Q����edʌ�
��.M����my�p���N�\q�?wQ9y׌��b��fW-�&�8�I���O���hL��X����3���`�3|���((U�b���JC���R�;�_��ﲠ�����H�RR;�ǻA��������
��T�Pf=^�Jʆ5��O���'��qt���%�9��������p�GJ��v��3c�,�&�����VnJ5z��@��u���N