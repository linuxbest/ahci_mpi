XlxV64EB    1686     8b0�q��ed�˺��=�ϽNt������،T!�]rV~��ۙ�.�|�
�n�[F���R��#暄I��q(�G�`�z�DC�e��_	��pxBU>R>b�xj2��Sn����ީ����c�c��O����K���%&VP����m�H]$��'$�[������^""��g^�$$�{U�jA+�����!�|�j0�k�ڨ�\pC��1����Z�X(������g��������Y�S2��lY�]����,�\0@�AA	�����p�1z:}�l4x�M�`�B��A��<��nԛk�����F��H/��'�K*?��qcq��Y�ڮz��QP���jkE'��*�Ӕ�}��+�uԿ<���W�SY���Q3�y�}5�f��F�Qo��c�4�i�&��]�B�<6Ge�o�O+���Iܚ���`vG-c7�ix�+��]�']T�Q2�hڙkљ�ՋQ?c�C|+�|����X����f����*z�����#���������6��"V ��_��m��ԃ�z�14��/�9��ݗ0i*7�d��x��NMb#��T=d�e��qLTk1.2��=����g�[�@w�%��� āT��#T���OV�p�?�s�!@��<7��W���ϝ�̬{�'��F�+�8��و+(���Lvg�[n~�.�K�#�C���;���ګI3��4�Ad���{0h<��)�N~@�˒ç�%�v��X������VPýik�[TԌ٠\����HN�N}����S��1�f�sA�a�Ɩ���鳕��9��r9DM�z���G��O�;��8��'o�j�.h_���F�S���V���b��żA��cj�64�yo����eBYWx���,�.ai�F�!/�=���s�	���� �u�иw*�����LB��XNS�G��կތ߰ �Y��f�uK9<�~F<ᯚ��_;5��Į3��u�X.!�!��c�j�T��㸢X�;{g��}���P-�@ST���d%�Y��e��!�O�D*(�|1���A>U�Sm���.�쉼���[��:s���'�V��L� �����eh�W�G
%3ޭ�����k�3cX�-t�q�B����V&�zu�vor?�N%X@�?5P�s���2�!���o�/TP:�P����.Ίɘ8	ۨ�!��-�+��J�Q��x��Ҥ���"�~#��!�웡v���R�@f����5���[��u�x�g�ԣ��:�w�RU3&b��(� a���N����bzzD��d��Q~i���^1V|�s�e@$w��\W�h�Mך#_]xm'���H'c��$zt��cV걪w�hwW�n�;u���JLYa�ɐ���l���ݿ�K�x	���F�Q �&�D�~q���|i:,7j�vz���|��i� W��"
P�- Uz�2m�U�q��A7(�r}e9&�kfߚ��V8 f��$�S��ضǠ#J2��B§d;��U4I���O��1#�nwl�4� 9��Q�o��z;���������u]�/z]�A�6��0l;9��Dj �
���Г��Q�[�j�g��|��`�]�4�Y�ntnc�$=���j���$ܯ-�ѝ�k��2��]�wk	�J�n��nԾ�y`)g	F�KJ*�c��ۅ׏��n�!��b���^������c�V�֭������FQ4ׯ�8m	�T��ADv�Q��R�(�=�c�Bf���r�z"飂��k���SQ��V}�>����O}D����6���K�DV��L�$���ݻ��%M)"�{�P{��|ۄ�
��K���������;y౓Q�ˊF�Q��aJϤ�F�G7
�{�:��so��0L�Y�?
��d}Y��t��� ���
C��'i���8�_!<�bU��鈄
Rޤ[_Q��m|�/�52�8���փ�MI.�[s��#KC{g����nf�8���Fb$H+��}6Tu����Լ�Հr�
,Sr��a�ky���l�:�A�����چ~sR�N�N�!���f�ZA��d�%��<�� �[}�� �^���:���Lj�YR�
 ��SK݌i�<t��Z�Q�Ϊ�xı��L�,<�4�c_����f��Z{ئ�)�+�{��m��v��g�ę
^{O�F؝[��{G!�I�(]�$)RP�W�߂RL���7L)��Ʋ9�;��	�Ԡ�[=�Ѫ~ ��'UC��V�`