XlxV64EB    5180    1220��0�Z�%��#�^�������2�����,^Ꝼ��8��]}%��/��*�0c���K*�>��֒~"���}�0������S�lĨ����w}��� ��<Ƨ��c�����9�<>�/N��:�i���?���(�B�[��&8�"���?E��~<0������4��:��mQ��(�B���ѫ�5�9qOXp�x=�ι��Hr�I�n�w�����-�ӏQ�.<��ybfdu8a���dy��
��8~�}s��A���n�x�oU�ͬ��HӴ������]���<�cY������CH��5Z G6s�pq	c_;�ԝKE�l�(mI���j[e�. D=!����T��6�����Kn˗��՘8v{N���G�2c��_���ы��V��hg�>&9v>�4��Goɖw�rND�V@�B!Ş����	�dR������]�I
������8��ç�	�|�KG�Z\�<�*�t���Ck��~%э9ә_I��G�P�H��.R&pQ�*Y�|��N���ץ�� ����$�/N��5�T`QۺX.�qs��(w}��)��x(u���I\�����K���3�b�^��sMRii.}W��5���9����u�5uV�-�'�ު��QM�Ջ�T�&���rN�����	��2�X6��Tk��'(nřp�P1^�E��1&>:n<k~�no������۬A�.%�"]|���a�!�O8b�)ʏ��%��#ْ6we1��]�[}f���WW�}VnH{��y�����.�Ii
��di���^~�����=Aɇ�`��gH�Jn���8��R�':]��lP��!i�t��`kyrGz�IZ��p��H0{Н�4(ʞw'��;bC���L��(�l��NSJ��o;��1���ɗ�`'�D2��˥oJ�{:F�H�x�;r(����u4�ew�6�b�(N��&*2Oɞs� ���P���^	#����(�H�'�b�-��>҅ȅ�r�rpIt���p�Ǟ�`��62m�C5~�G�L7��,C�k�L��J ݢ:�DQ��Db:T���rb�3�Gd�LO+�Q��>'��<��+~,��JP�� ��C�Ѐ�BY��"[�������r�UUG�E,������ï\#��]��xr|�|�j�����hXX�$;�o�iz��]�a&�,a�i����]�h�S ����q��#�Ψ��]�g:��HKcQ�ib��ְY���ݤT�{RF�Sy�x]�a�7 T�Nԡ�|1dMl/����i,M�'$%]������]�G���W�"���z�$���Bܖ.`�`>D%/�ΟmL[jm����hH�HM��J��v��t1r^#���mX=�|dh�3Q6�����}�yNd��h���C��4�P���L��~0ou�J�g�{��́�a�� l�m]h���~�� >�d���B7}�:'9�M+��hQՑX�X��P�6[ـ��kV ��)I�܅�)�׬�f[��Wb�%5hDª�f[��jI���]��l��r-�=��`��S��N������IH̓�#B��21�uO��M���z[��Tq��<R�1�3w�{�|D�nŲl��~w��Rf�g4rs��Q�.[����ԫ��\�]/�M9I!H��-D��hX�C�P�6b����6���b��q3� nSS��I���c'r��:�e1cyY2J�L@W�O��-j��l希��������M&F�IT��H��ͦ������a���Of��b�35�?��>D���3	�i�3�9)@Š��V*K䐮&,�<걥� C�ݤg�2���78t��2?��acδ.dK��Ȗ��S��Q��8<��w�XХ8�b~i/F{_7(U2̏�s�ϊ,R���?
����>e~�M�3gm�@'5����u�sr���O�cI���f��1��d��?ʳO����*�̕�_t�<��2J�Ƞ(��#�qS:��{�A�@ʄ��>-J`�jCٕ��4�
O�H6�d��
�z�.�ֻ<%M�j6�q�8J�C�Rw�2��ALK�)*��<)�@;�-�	�	+ϼ�3X�r��3Б��l���fy(7���^W�a6�qMr-]�C��d~CR��B3��z���\��#�[�<�Bԃ|oz&[��{GX��c��+����e��o�A1�d�Xh
P���~mÏ��]-ۄ��r�L��{��L�:
qW����oe�����0.E�ǜ<FZϓ��:�&��#�m�r��H) �	�����_��$O�cov)6C���j
���حbN�s�dmM�+C��$���t�������EG�a��������:�VP��:=�����)"��XYB�t�_Eݟ@#F{�u��"�+��ү���)S���!�a9Ҽ&�ɖЖ+P!e�Ca��'g{��1%7S��7g��v��*^67Z94��Ao�@�eA0�	�Q�̖��=x�=��I���v=����֌�Ȝ+)��ת�Ú~�5�ʫxZ���ѭɍO������γYo������A�vіEL��.�����<�ΰzuc]w����]�t�R�?tb�v���3G���>?�o�#@M�3"�Kku���G#D�HK�(�o^�tQ��"Il��Rd5�{���d��הb�7�YMZ�<����֐����_M�Α�uٚ?!\��ƞ.=˼���L��q�+U'~\�K��[�����j��jwxl��B�8�L��Qݻ�<�f0�x����{�����މ&C,�{I�~��JL'���H$(E�ߴd19-�kgRGp�}�L}댝�CְA�'�(�p7mIr��*~u�� 㭄8p��m�g�����v����e�OX]�Ɯ�u�\ܧچ���ɎW��r�W�41�\
��k¦
��p�W���*8M��z�!����X�رP��ТB�a���X��JI��j��F���b�Q�4lF3d�i��ѵ�x#"/w��4v�G�ܼ�K^���?������lL�
�=���� Z�$F�T�巋C,�
+��G����0���k�_�~<�Q֭t�����P������Lo>��\M{�]HAM�+�1|?
F��@L��M ��ٵ�VЄE�)�}I�X����'x?�L�Z{��$p*�P:��ڋ����
"�ؒ�L��(x�X��SN/p{D��S9�]E����P4�d��ϳ��6���j�2(���G���q4� ���Kמ̧�W�7oX{��mG~E�=�O'��c�*��!JP�:$hb{�J>�G�jΫo�;'D��n�Fx��bVԊx*V��ʱ�w�P��d94�<���hA�����F�D�T*�9�a&f=u0Ƕ=����Bqj*0��Č��}C	Uu��q*O����D��Or���a ��^�G� o0�BZd��*�6M�p>�&L,Xzs5��g�2;�ӓ�ʟg=�����.��%�1�*#b	oZF}̑txX2٣�V���Z� �=ϸ�a'e�Zg8��Y��S� � �˰8d�U�LE'	�I:Q��RTz�A���@���z��SR���QҤ}J�>�R���Gj ��"#�q2���]6>Rq��� K_5b1����3���*� 1
�, 1F����*��`˵�fāX�
s�6hd���lQOh�*v����w��-,�	�ච�d����$�4Y�Gr��Y3��R���
 Z�Ó�����f��S❿�\����k������t�".e~���m���QEO|O�z�y��$�?0(�td��7[��?���3�EjDM�3�F���S(��X��dO�j�����L=j�O�r��}�f�G�I�>�qZh@�{}Y��k�10�	�BLM�/_k�}ݢ�$�	��j�4Cc���j�b�MҊ��	=���s՗��H^��{�"�_�C0�>l�5��֤>a.���{.v��_�eXpD�^(H?_�L8X
����`u��j�gj�9�	 ��[������|� _����Krf ; ˃�b�k�<��I�V�Gy�<T����<��<h��[Gв�`�z��R�,��q�Q<�8��s�/EE���hyYj�F�`y;�%�Z4q���F��X�F��[�"�֜��`7%��;/}���C���;�O�C�J���59������Ek�Y)W��O�7'���E��'Ż�KƆ�g�_�l���a��m�SF@k!1>@����}��.���@fHʲ~\ ��
�E�.m��	�]9'hI�q.$5d�i�PcA�pB�t��H��	��y����Z�',늢'�rԡ�r��p����9�s���]�e���向�@��]{?q��ʦ��������2��f,w<g�n��h�ڃ��Ku�'��񉷗Q ��h�}9�>�m��;��O�M>��X^�n�Ǹ%���2<�x�-&��H�,n���/C�z����+Q��z�\�����Ȩ������d�&p�q�]�K'[8���'��Q8Fq�y֎6"��i��Oi��`�b���J�����L	��폯�X��<<��ф��2��=�