XlxV64EB    156e     860S�kGu7�P�R}�����Y�~ۡD>�YN���DNWlJ6-�PNw�� a�@�ߤ���;�4)��z�9j�@h��w̥\~��L>�'Q�����`�%���� �����C�e�.|駘����X��25s�P�yP x��
��=�:���I��4z�7ݳ��h�#-a��6l#Tsk�������O� e�L�IU4������dWפ�{jЗă�{z� �gv���ws�#� �s��l]���Fv��H��2"U7Q^��^��Z4�DN4�h����HDZ �H�2%:�A^.k�&���;N��c��ǂ�MY��vZK
p�`����gZ�d^ä?\�\�����o}��/ ��$�H5mJ��7�4?l��f���}��w���X)X�0��Xt%/�r;�Q{�4P���!�%q�s^������i9��+%��x�S?�������T�F������~��Cop�U7���I���nݚh�a6Ɏ�`�c��T[k �I�RI:������%Z��LDBl5_tV�:��X'�mD�c�<�.[�d�9`�:A���_5�ZV�y�������'�<���KF_��*8��1�+do!4��-�n#���_f%�
�����-Ōhu}�l�:�ʤy�7������.bK>o�؉�_Y����u�����;ªki�,�z���{O �_�Bp,V`U�8�]��rl/<��w�G}[�p��Y3�&�N>m'�0����Q�Ho-��>��=x���d���D�.�聯����2d��'�JOv��7��jo�[�~O�9`�]�I.x��U�����J�,Ӏ"i~@�(��W�)�-^ue}�.79��NwEʽ����=�6�&�ខ ��]�<<]?�����R�ÄQ���D�B�INs������|Kb�td`�]��ĵ[͚���l��Z1C�r?��C�M>�)�[����"L��0�RW&Y`����Z	T��d�Rg���A~����w��� �� ]Tv.�}o3�~�ã3qj9&IyQ\^�� L٫��X�/�&��k��I�ˬ����m������4�z���0�g4�%��@� ]G�t����ܽ��q������bg�b=`�$��~*��ʲ���|	@J��
�ʔ�:;s~QcQCYzB�{V�E��%����!�<�BG�h1D�<IΒ~��ToV��<m�Z�	����^�J�5�7���o!<M���J�G�1��:
��2�[���o�g�L��o[��6l��:Z�X�[&EUf�"K�q�Z/����9�	�5]T5�:1X��q�i�������N�����u���2����bjJq-�>�ǝ'�{P��s��L��5Љj6�I�?��p^t���=��~p��v�����_-K��*����jS���3�z��~ ��CŬ�.����}Dz��!x�
��n�PM$8�s�Z��=~(��r 
���i��X��Ȧصpe� �
#[���؊�Q�P}�i�<��Q:/��	~��xxi��v|�x"�	��wh��.W�\c\�<*'�) ?����M��4�|hrZq)5 _�, H��-���Ј5���[=���z;7�|.s8n]��u$� ��*��X/$mr��/:���!R��0]_��R"�R�؂���8�J4��	�KC�=�o������<����νE�+�my��-E�V`/�1N�����^���U�I����2��5ǎ���,��������(V�)Ix[u�`��7ƒ&��~�>{��AN�����$��"6S�i�=�^P���n��N�!3y�����!W���H84�E�0�1�O~&Su�>�8�K6<��)1)�?�/�d���'����V���<o��l�`yVicqE~�d�z�-�����+�b�>�_-{�������r�����F������?���pI��k��AiRlʜC'%Bs{k5��!���V�o�n;��������RU��ȧLav�ɺ�����,n�pÈ��e�v�(�Z�5�zqd��3�Ƿ��2W��Y�9��Ke�o	AP�[��^1ڕJ��O�A�I�H�7/Nr-�'�'Z��8{'��e,�{ƣ�