XlxV64EB    2832     cd0�T�~���2u����N���1@I�jm��<S� ���9�U*�~ �@#�j=Ɛ���yt�~��$K��$��2G�"��K�<����|�;_Jd��=aE���`�ɚ~�ҿ��C��P�D?`ns��s"�*��x:�F�k�l[�Ko����'g�9�U,��:$sDPN:D;�=�ͭ���[t̜�w
MUS�I��i4�f*�`i�|{K�<j�Iu�U��6���|k�*Z\hm���a4(W|��NdL��k4�r�v�5�X�(U�1��я`O��2N��[�q-���L����ި�ħ���ޖ����n&��(�<�����?���w���qG��z�'#�K*zN;?d6��$��C<��g:����o�L>t�a�D eB�z�W5�q���W�|
*?Kpޘ6�T��z��W�D�� �9�3a����P�H��"�λS�=n�Zr���@�V跠�UY�:11Fl��*Q�~��f✺\�����!iƊ@�|t`�m���ק����P�<hZ׵����u���ӡ�j�>t�d���i�_�BW +�n��.��8�CG\�>r>r�\�T͈�c��s��I��2-�;���5�B�+�!�M��=��pp�<+gD�g�R�	Db��&n(�=7^�Z"��~z��X�� �W�؉�w�}>(��"�-���]^:>�j�k��SYM'�-��{����^�Rf��y7�ѡ���`ܜ��<�������lE�I�Ń�A)-�y4��Y9ʾ������(������ڤ ���g�){���<UQԺ�,��vq����!�E@)ə|��������~g}�f�����٨Ŝ9�q�
)��E*�DM�Ao\��9��m�o�U���	4��l�	�n�������alZ���A�`�&��C�pF?�����Uކ�H�f����)�>��t�uS�Z��gS�a<��L�04��n��6I�t�=�(�-g3�&(sc�;H��ם�Y�����T�G��~����� ��[ie�4�w��ݥ����ˮh�%�9�������,��$ʃ{���y���^N4i�a����`��3����[�rC<��J�nV�|��5��ѦY�bJ�o��~tj^B(���\�]:IiĮ~O�ւ	Y*ዮ��R~tA^Q������iQ��	uC��r�f�ol�mr!4>��� {[j�8��[:����:�yv,�,(`�����S3B`4ѡ�܋���ʃ��Ƃ��v�;`-�BM��m��������D�?<���GKϺ!}Bp�߿�O,E�ْ���/9:5���w�>�~)����M��73
�
����<�ȥ�[^fA���e�z�w$�N�1Aum7��늄��7˜�oVT�����*~D��?L7��@��"��(��M<ȍG앱��T�� �n�n�~��݊��
݌!l��_34�{�'Q���D<<ƹ}Rq|�@`�x@"���Vj��c��XZ��L�~��lv�~f{���yO���Dl�����t��0�)ߺ,���[���ŗ��������g�s�)x�FIŒ2NZ���b�k�E����A	�TO�j����g�͗�!��ao7xᩆh�!aZ
M�=��W�˶:CK��3 �49G���)eH����F/�����]�9"l�B����{��.�4}��`c?�R��m�����Z�o����u0�
��0��h ���_�zv���=�!3P�ހkD�y�|������s5_��ϢLH�+b;��Z0�6E�ԍЛ�n�D@ �/���̉E�-���I���x��\Ih��5�OJ��>�0N���d�|�r�'_�<�>��fSH����1�}cN�*k�I���2A��ϫ�����5�rj�W�K�����\��7�qd#`����U�pn���O?�J��[�I�e5�湆���͌�!ʔs����)��=�@��슩��eM��"�]Rh�����ro�#���@P�m�|.��1
��q��p�'�Sԑ��k�
Gw����,�=E��N���X������4js~����<J�wSC����~ʇ�]I�����L/6R
��КC�4�(&is _V(DY4Hu
�RHȫŏ��MQ���W�:e���.�e�RO���G��]��:uÑHd��NV�p���Y�X00�i����LdMIq��}x=ؾ�w3*���Zq�t��]jky?�:�ҳ��d�M�u�vȞ���P�\�:�����u�&��Z����$�*�8'75h��θd�>Q��b��%ۊy+1��/���
�c�� ����D�{1;ʠ�b���Zc���:K����O11�e=/؜����H�̘RTOٝ[� (YK����p3mE]������]PݴU,MZ3's\�@"�-��U53o��Kl\�%��Rrw�8�S�&�0���CN�l*�P�K�v��p|W_�����Q�����Yf�9"�O�� P�K�Xꚗ����1 m{ݺW��ϾJ=%��%�'��	$�Ÿ�ݮ� J��v�Ú���F��5~�R�^�-!�1��Ň�����<����P��KJUmc:y�6���>{��������Ԍ���i{�"�M�"T���za��dL"?-���(s��?ZnBaFI�v����,�R6�F��{�H^=����q�b�6�*�Ϙ.�o]Pd����#���	���̀SU�1?�:(���aL+H�w,�d��gڑwBeB�d/����k�":���2� �Ώ+��"�n��)|g���z�̾��)l��9�t@��9�y@:	�
�qU��|ȣ����o<%����;l��f,߳5FŹ�,���C�8H��23<���9��j�S�3��y�Q�>�ɚ����P'_k��0�`��(J� 9�4����(���Χd�����I���,���1��B�[)"�mS�ݳ,4����{�S��S%��e5�3	 �0��b	��
�S�����t�D�D2Y��\�
�݇	<�N��JE���ڡ�{k<�bjF���\V����9���@�Q^8�w�FMv2��`�?q��ۗ�e��MqvL�
g\,��%�y�8��?�&"?Z];����Q��Y-{d6	����β�'��<���
�������$�Zȁ��5>�8�7Ig��lwB�;������_��5	R��5��8�C������=1i5�)+@�:���!1s�.��V�`�0b�����4T�
���QU��>}R�5u��-/L