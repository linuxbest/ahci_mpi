XlxV64EB    1d25     9f0�_���-���s��y�L�\�bH��B+g6����C	>Q�=t��^�ф�ǈ��]�0t��{?��jR��ZD���x0��f�}j9�����;ұ#����i%���ʆw�4j�ߛ�ڟV^�sڍ�V����+ޑ��
ٖHmX#M��Mr��\�ՇOr �?BhL��\0��#  '�]�<+�w��������3�o�,v�G�"��oz&�(;��u-�a�����@*����S��F=����㦀�'}:
�Q�	r^������-�/T� l.���'����yNܸ�^�Y:��,�2�zu�:��~j�J��S ��|X��.���?x�D��`���4���ݛ����H�fw}��Y��k���l0"?�j���r�Ժ������ƚ�]%�����%P�b�ߢ��k��ڀ�'!����Ufrh��D�'q88�H89Q9	צa�"���$<�W��̂z��`�����<�d,E|��E���I	�ߍ��{�n�jջN���EcH�;r�a��['�M�/���w����4'��O�y+����г&��:����_��!�����!A�@�?�~ud,�j
~7�j3d4���;�O�d̽OQ���R&����ܞ�hb��
K���BB�Y4վźx�,�Gn�/��^	]cӓK� �Y׌��I���9�B��x��{k�+#��!���{���������K��NO!�q�(׭k��hc^���<J�����\��	�@����̚���&�3}g!#n*�9��{�BE��$����Fx�	Ԁ����'ۨ0(��jXG�T��b�`����q��&�O���J�+��5�0�O�g"j�#NvS��ɧ�N$�y94c>�^�.m����j�̳; 2gmj���x��S82o!�E6����i]��^�4��=x��cԲ%]���'0�����Ŏh��� ީ�Oʟ�'.2D�A�uh	,#�\>��)k'�x/2 �=��$3Vǹ���͜�ɷ e����=\�%}�mm����26�@��@����M�$��p�O�'���{���f���ؑ����z�@D��������W<}o ��E �xᘻ8s�>�T���\?�b�1����6p�-��i�-��kDpd�dƸ�d9d_�jg+bg2Y�!i��d���wg��~޳TkN����A�	����o`mR0�D\z�xȄ7��H
(�Y�Q}:��)��)��ݰ�]`M�3�\�`Ĭ�w�3H�~I�=Gءft��RYzf�ϴ7Eȸ�"���&�!_r&�n[�v?�\�f�đJ�����D\�fyt�7M�|Վ�?@"Q[��Q�<��@���H{8�F	��}[���V Ћ^q�͏���6P����J��(�V�*�o?�\L��� 1(V�	D�����R�8*� N��-�tx�h*al������.�uM!ŉV��ᠷF;qM�]�|(g>Z`"]M
�]�,8&g��`Z[Hb4pE3.@2�aUеxN����*r��-��4a�x ui*�Fz����� rd��}�.�V��3����v�Gg�����z���2��������X�ARbi&��\u�⯄����˥ݳ\!x�h��v�$��ĳ'y@���ov� v�6�g�Fl����4��0�Zp�#�:���e�����0Bo�y���F
fYz�g�p[��bGE�A��b�ue��O������t����-���h�J�V��o�Z��|kI�����/g.���E$��Cy��٪�f�:�|���$�,w!��zU�[Y�E��ި�Qs��0 0�ԊY����8�
��u���xK��βx���Dsm䡡B\�ya�DP�P���>s�yǃ-|J!.��t�V������z�^�<̂��78(n�Eg�"	��`�':b��n����0���a�E�A�W�V��E7&��B�zO���l)LZ�m�}B���'VO���j>�H�a� vN'�B8^�z���[��jɒ�����g�������6|0�&���5i3m*���~���������"��&���x�~�����J����/��ݹ�A� ��Ȇ$����&�o�z��NH֓�˻����b�����|��v��.�a���p�ݬA̖a�M�ő)P�b%��&��-������bN��G�v�m�.�g.�iZ�N�9�P>��/Q�pQ���b�%�}!����pܡ3$�K����Q��y��ѣP�O@�[�n���8ɪ��C �n5���O�o��,I��J<���(�Sm�n����H��a������W�n�م�n��E�x�
�,JM��lT��Q���f-��*K`����U�4B,�^���b��t�%�؆W�����V���&�B�\�J��~s@���e��Ȇ�i ��A��� ����G�̨?�Kk;���'��{S�(���6��@�2XhYn�p��W~�o��9)ނ��+�˵�Χ�2l1N�ѓ��J�P%2�GV�f���R��,Z��u