XlxV64EB    1820     990�+~E�@��l�B�bt ��Æ�������� ��L_V��F�M�X�7p��\F�K���bG�4;ϿG�p^��;�y�s��_��F7[_���No	�|�G��F�>v��_��{O�H�+w�N�+�-�Ũ����k]M�Jn��,�f5N�y˴˓�%
��Tx�E0���R�xOK�RO�3������3C�������OM`�Hw����M�]���zH1�`�r/l�� ������?���Vү3#� �y]��YF��M_���Z�����������i�P�$�5�����B���?�HqY�*�b�&���ݲݟeᴽ�	Nt���d!���\k�-$�H�'3))��
+���d���Pp�Kr�&�'�M�,w!��𭿄�^!��?�+�,V v�MajG�W�e/�7;r�n�$�Ɉ�'~�mY�(�E�����,a���\`L�h� =.�V^u�kC������h����;I��hm.��l��Tz����L��C��B]��$�{�0)����uܦ��6�e����v���VJ�� 3�1�h�oV�K�a�}w�m�2^�E��1��>�F���W���� x��%;eW��߿�j���z��N���o DP�����"�������x�M�I�N��Y�l?D��ٮ͠��U��CBꪹ�a;�å�Ơ'Z��t��'����y-lG��f3A�'�.d'�XQ!\\O;���2��B�2�蕝u1`IF
%�����V:���ӜcS%�q��,~.X3m�wc�J�&��|�o{Q��拉wۯ-�:]Ĭ��S�5��P��}�%A�$�~���J�/)0�:�I���ªq��P3�_)��_v@c2��vM��|Deo���i�%��D���f%D��oj��9n>4-ھA�eɗ���&���l,m\�R�Uˣ��o�����z]������,�\PhL^���J���=��#�Y,ħȻ�<a1�ϥ	��D�i�,~���+� ����tP_���k:�2cv�Ì2��p�z���$4��s�l�o'�\pe;^��V�)]B'%��@�C8��Id0%��u�_o��둰X�jx��`����6��c* ���n�л���R���h@�mznzB�k����ݘ�+3�A�6�\�(��mA�]#��U2����v�ma.�?�?d�6|둖6{Jۀ$�������U58z�-��@_��A�%�-�In�$�1���R���6i}	�cg%}�7��cJP�_ǘ�[�ɗLU�ׄ��C1a�|ܪJj5�c����
Rkq",�!���Z�R�ʞO21Ž�F!a�D[��8��1�!m�KDp-n�� �!J����b�v-�ST#f���Ž�j?�Mƚy2)l@�=,��nq�r�5,��h�0�_�]�E��{�����9`��-�Y�缋^�׌��M0QTnd[I�_jmlI��[Jg�ie��4wY"X`��򭦉C�CN�rդ��A����I"�¥�SH6t��\�.�Vp5�~w)��F��-Yn�(T&�lT�0��4���m��?��p��+���_[�ʃu��FV4�n�V)�٥lst�:m�=]��<m8?/ڑ�'��Q��"�
��f����O�`�l2;Oiw����u�k�~$��\�>�,	1������<��.T�f+�/B��޶IF��� �N2��Ř����\	-FQ�zж/��^N�� ��L����ΝC�Wh�v;ʃ��J�-�p�^6�&�|�0�N��٫q�.PanR	�I��H:�n?7�a=T�rY����<A���4��ϳ'�!NQF�cԖ&�X=��	F{��yn|V��ћj$��TM�}4S�Z@�Dk��!_�;k��{$�]�,"�3u�.H�*n���J�7[��X;���I]��O���4��E��a:��rY��,�JqQ�!����OBT-z(%�"��i������v|wy�.P�7��
�p@U�(rDC�n0�z��0��R��b�����)D��1_4�כv�W ]f4�^z�}%����A@	��/u0[-ò}�0�S4�Sc���hfLF��@T�J-QW��n�Fڵ��ѿ�� �,�F%53��h�m$�W�΂
�M$�j��Ҥ�4��WDK���W�����ƊE�8
�Y-�y�����xf?.=��N�~a#ОՒ�ѐ�ϖj@c���|��J�PƑ0�Mr���C�H�� �#���b���E~��$8|��S��%tES=|��C�c ?ɝ����q
R���T͓�����i���l~Y#��h��|�ܣ6Y��$�}U�jM��g/;�P9�X
�uo����7�v�P�������j9?��� D�?6�R�㾍��Zjh�oN�:ia���6W7
� ��;vݐ