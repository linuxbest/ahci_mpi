XlxV64EB    159a     840��JZ�B{�h�0������h��'9��$��h�:I�<����O�de��&X�n��#*��xZI,�\f��a�Ԩ{�ziТՈ$����c���^��GNm�eȃ�u"��<ѐ���������p��椓v%�����zG���C��6&
��B୾��Р?�)����]�\[���V���1���܄ �_>lS������Y�)<��4R�4@��zg,VK�V����G7K�|_
9���j�VKC�_nj�=��-�q�6��	L���&���b�j���8�,ɇp���ANY2���L���l��/�7��S��D�#�Z/��%&�F�+_��)j�<�C��p0�\z�y%�U�W���$����H��f�	7i��.�z�[��ݥq׼p�HFQ%~+c�3
�y�n7aQp>o�奲%=U���EG�ps�-�!t��K�$K�:��%>�Mm��cXNp�q����W<�\~y�zBy���)���r1l�n���r���u&���������j�<�L�T�p5�y�G����1 �Ƹ@6__�r��D��N�H��6�l� h���v��ҿ�I[��8c
�V�z�[5�o�v��$����,��eD�P��s���.�#���I>N�9w7xSo#˥o<�}rV�6:���R���R�)�`�?�0�h�p�N�*�;/٧�%Aی��e�J;����uuu�5�2��PRt��=�I�c��ħ�A�q��ְ�|$N�����tޯ�!���cK�%)"�*�l���B�ƀ��[���b���H�c���͉���|^���4��/ZJ�ğEp���Φ��գX���Ċ���W1)>}��7e'EŢ	��ܠ�����8��n]��;��Tέ>�)T���99���F������s��V��Z�Z�ׂcC#m��0���'�;��i��vQO���=�֝=��J߶�'��(v�3=�z?a��T�E�TR��v��f��Q�3;�C`iJ
p�uQ��hAZӼB���$ӟȿ�v�!����BV_A����7f[5s��s��{�4ȄE�6���+��Xo��-�C��V�ioζ;� 5��]#��?!L���b��0�j�}1��{�g]T)�L�)�M�8U��=�n�U�Y��l�"��7Ӄ�XfJ��	{{}�""�$��?O�5��Ꮣ1���6��FC��ו�V D����Xw�b �r���]e��.�sP�ĕy{���B�ǥ�d��[U��\,��KƏ� ���V�H�q%�?�T���,C|�rP���)�^�X ��t�\��E<�sb�ΗH�ό��]G�{N�hpY����t�bQ�<<P?�Z˭�����@���T�t~:G�b-��eV �R�a.וÓV�=q�#0���k>�	�u��!���3������i��*,+޸<�gw:��S�p���N^6�R8K���y���so�q�>ل|�D�.Ȏ3ߑ45U�M)���Z[�DW)?��Z���A�og%`��1� 0O�\z���"�\Ѱ��%�����8$g���^�{�py��\ǋ�!�[�y��'�G�H�n�Q�|�rr	���9����N��^�>���Q~���i��ߩ������M�5b��"�ڹ�����������)!i�.�d.̿\�zo:*�&kz*��!jM"���C���E�����|'W�ϼ����^ꗨ�:�RKo��f�k@�\��$�{��uƊ��Tc<�'�.�Y��v���K�\��/�������2
�u��P�+�d�@эY:��~7l�R"
߱~���igj[cD��ܳ���X�$��H�k����Z;Ҏ53�=�sh�(�e
^l�ӁXw��C�,�����ɧق�1���Dc��#����P(in�4�_ÉW�"�t��ޖ�T�c�B��lo�"��g��?$�	J�X�ԎX��N$�1<�|f�����sPY·FM>���V>1]�[2x�`��`�Z�Ks���?>�_�[$2�S��$�K��d��Ug�N��mh ��`н��M�UE8�������0�"��(Ow���O�%O�dt��p�٧vY)U�j)F��ύJ���