XlxV64EB    2a43     c30yu�d� ��E�Pw�Ew��{ua��3��P|�4�2`��� )��Ë�H���r�<�k�&�a1�H��[�`��\�ǘ���:$ɺ�g�T���a���g��yaIJ��&"�3�~����f	���v�,�±#x��5A�t�������\���/��jch�j�ټv�qlO(J�R�(L����
�m����,X�9&�X�uu�L�֚#ϯ��×��ί7&�c �k����݌�&!U@E���F��7 �~��Y�+J�����A��v{X'`jxmR�!�(��w\=���G��6���еJ�ѩxy]ʦ�kM�V��:����"����Ѣ��qLU�A9�O
nVI�88�)�h���n�9xٚ��}	��>Kf±B%�F` �&8�~fn�7@"(�O�N��W�V����R�j��7�!�1y��4iJ������G��g�j����N! � ���<����%,�����pL�~-�����Y/G��Hm�m��sT���v��,��m7���x,�'�=p����e�;��cbw$]%X`�,2�^]�z�Q�N>�M�E�e1 e�ߺ��f_��D5�H��ʌ��`���˺4$���G-R�1L�ϵ3'ǁ����g#s���,i�o=3�6�>���6i�uFKw��sN|���q���`���mp��|V-��9�@�����r-M=*�݇p9��~�+�$�2Q�K����[��"5C"X��T-J�_t�3�5�� �l�hGۙg?`5��}¥�ݗ�aE��2��Y �w$���SC�L[��D����P��m�I���`=śYp\�-���%�u��m	'���-Z��`A!T���Ĥn�"ǚڕ�ߕ`��o2�
�6`.࡮0�E�%,XJ��2���d'
���b�o����|V��|�.'��s��N�|D�6v�D�~ο�<&�X$Lb2 �Hoj,Ne���#!qK��
�Ǽ�yT�f��^#m�|>
�̷�`r��FMƁ�Q��W�5��7�	
����3l�������o!��6zJ�$�Q�p	����(�-Si���3�� ����]��g�l�@�!0<3%��ѿU"Dֺ�Q����wWi��6)Y�
=/@���v�(~�r���@ef��y�q�P��I<�ӷKzß%9(�����QSK;�]J4zg���Nz��x�
���4��`1�u�i*2=�.Ǜh.A����_xFj�(���B$+�"GG<#���wϗnP-i��*6d��]�(O񌞰���	j|���?��d�q�V�7��t��B�Bٗc��NBQ�� �l�y".����捴�8,%<?�d�xٷA�������ݪ���ᔃl�E�K�F�B��������g�w2�=�����p��緓�e���ڏ�D�����ʧx��&JRXQ�����op���$ʾ����M�1��o�|m�[΢��c9�������8�Q�J��6V�@�{28�
�vx0���.��p�3��kx��}��vWt�2D�ڒ��X1Gv���	w ��\ѢZ:����"Շu�H3!��a�8�]��7���'P�:6�o�n\�Bb!e�E�nB�`\]{�YAx0Y�ȹFq�ٛL���`�a��?��
�D�5��0>}���8.����~JMt���ʹ��Rf�+��� ���WZ��3���6c5wB��D9z�e['�		|l�JO��3dJ��z�Wz}�&ny�A'��}r�U�E~��I��5��2�QN&_�r����Ӯ�8�7��*�\se�X�Y����AB"�`81�ڑ��%!��*�T���C��k��V�����3��:˧d2ﮤAgO3�4˔�I�� yЗI��>�*���F�-����G����L��t���;CBoM�Uf��a��0m7D��f���[���k��W�τ��6��xGݤ���"��_^hMU$cU��<�QǏ۠��)�����Y�)�a�k� U��7�e[@���I~	��O��&��')ڴ����k
�i��ÐM��+��.7U����D*��a9:�%���mS_�ί��v��P�����?B%6[a��b�ݚN�y�`w�&|d��ir������j�RU��͘S7��Z(��d���ؑ0<����t�mpxe�8DJߑ��~���7�Eͽ�n5�fC0�z�H  ���"3^��ry��م����T��8�U�V9}�P/���t^���ԭGh��k�r�e���C
x.���)���`�l(?�Y��+�ƚ�ߢ�v	�욳����ٿ��m1P6.�����	�\��Ok�Qr�����X�`kb%鹫�� ��~'n���-���+�V��@��nʚ��~���!������n��\EG�p���=���J��*��e���0���=Tc8�0k�e2(��r�}�R9�lOވ��m�:)d2��1S�����Z��1��P�QԾ�@�0�m�z��<cS��/���Z�! ։��M��wʖ3Wg�1���/\m�KS�O��X�`O)�P��5	�Vm3;�N�X9m��s��H�o&aS�#����{�̣�&�`�K�W^�4h>L)r��p,�~����Ku��Cɷ�r��*�_l_Jw��(eil5��>��e戀8׫v��`QJ�|�N�]�|���CJ�<bd�t��� �8D�5R������H�\X�������<��|(�&7�z���"{�*C'�WW8��au>�:[�÷�dI��D�Ld���7���9)3~��&�����sQҵj�N��DD܂eg� ��3�"�0�b�Z�@`��������0W%�hT �vm3g�Ips>s��N��\Kp�aA?``����K5=4��b���:v#��+����FP� �[��X��p5����������Ѵ�g��;+\+�uf�or��8��*��J�ЪJu��fK��0�)��#F���5��.�uXpq\%�����Lܵ��/dx!}p?gE���v �1�g,[��T��FuBi�O-�2g�=xZ�2$��ƣ:M`�Nw�N&,��խVC8��G2�(6������z<N�ߜƳ-�/;z�V;