XlxV64EB    1876     8e0^?�B�eecE7�,j��~,����C����<Ct��sD�=$My���ZN�xu�8؃���s+F�:�P��A_v�&��Z�TE��X�������[>�E��<aW�0;�����Q\3ZrlG;��tjt�2��r�E;j�U����I!k�s~���~�Ҡ{�r�ו����O��j��X����y��qZ��ۇ!W8���.K_0�7���Ue��l�$� ���F���1��g���\X���@C����U�#V�Q͊�۩�n[`�îk㦥��,����[��֯���Xӈ�����M�woS�i����`�\�m��?���Q�ї���]�F�W��	qq|����1̫#~Z�_E��u���c8j���Z«>$%EsB�Ή�F"4����wO�/}ˮ �̖��F�z�B�}�>j�w���1$��7���0Mb�uWRM��^)޿�
z�lI1�,i��tq��z��������uq��$(HG����rz��F�ͬ�t�9��+�E8h�1֚}q<�N���$�غxɫG�~�{��οl��| +޻z%�����m�ڔE-�YLjg�;��9oFrԤ=�?�3+�Hʣ�Xd�g�!�BM�t�8��>s�8��NX�����H�������G[�{tRORn'x�`lI;/�-"�?��'��OMg���|?�N�� s����]�5p��MsQ��^,gN�ܒY�i�b.4�X��i>m�d��>"Xp�m�܌�\`�ձ�`��;�6g�si	�b.�~�	���Ҏ�O�C
��Q �v�YY�����B�y��PX����C.��|ʀ�`p�6��E"/[�u$�7���|�S�:�O[o�Ю�H�Y@�P#c��C:�:#Ɂ�S�!���u?��d�+�town4��cD�������
��	��Nj� Mצ��GC�y�1.57���2�ϧ0�ic�'����jo� nA/�.�13g����:�9����&ȣ�0��yL	��$�h�
S�����gŬ
"���T�W�h���oB{ii�%�i"r`�$�T��P�P����'�����J"����V`���ZO�ֹj��ڧ��/�7��	b^���A*5wݾ��E�R֮L����	c-�PQL	j{S!%W8�l�O��42ri
:�=���娩9�,K`auݖA��h��<徿���`n�(���M��ڕu����9��P짷�H{!�t�t��lP���lP6�vݶ�����D�8v;�hkx������eFeW���Z��n�'�c��O���n��*�P�n<�Z,O�/s�������tS�纟`6��uM�i�V�2�A���o���'vՒH�`PWt �� x�S��3Zܜ�"S!`�:9k�e)���XR��t�ʓ��qk2W���J�h��R�8��m���$`������8aȺ��@�.����?(����ج��L�:/�7���(�~Gf>�Q�Ĥ�N4r�����k����7!��"w�:Up�T�J9�O�/���m�b�s:�����w�ϲB�Ȳ���k�U�rG�Tѐ�l
���f=W X-MٽJ\��⿾|yc0���|��Z��
[�5@ퟑ��iRtdJ�r�ل��#_�J�D�z��M|@���`�ƽ�=#@����h�7:S�:Ԥ\��ጒ�SU�z�/�ȇ}nU�ج�	��nhd��5^ۍ�Zz� fTmo� +��F��()/�-�<M~F��%����"�"��(J�d����i�|��oHG��1��޿C]ݦ��R���y�`�R���	��]��	�Q�9r�|���N��Lu��f��t�����Vy��>��{k��6��x�#ә[`�E�SK;��d�n�xԞ�4���5�=P��:�<*�D�b�k�����o�[r�(��� n��1�QJ��d��G"��3(���ZF9icIY���y��E[�gMD�1�s�L4�	�3i(������mqy�H�1ۺx+��)�0���Y����O�:��x%�'D�Kn+	X� =>��"$-փ��
 @�Zt��'k���x���bb��亟��m��Ԝ�P|X�ŗV�����r)�ۊ�K�E�=ĝ�@����p�a�� /&Ϻ��^#��;:��2�W���%�Q�����shM�^���:l,w��-���n�5��w�R��nŇ�\�/[f��B�� Pcʦw��"