XlxV64EB    194a     9c0%����~�n�D�*��\o�]���J+"�Lԫ�����;j��2l&�� �T��OH7u�9߀&�	�g��77ڰV���{vF$lm�N�\�}-d[�j�j��+0v�\>�ʣ�W����]�ð>���d�J~�(+�cUmy�fI7���P^�2F]�ĝ.�^�]�5�ѕ��=�@�~�#&�j�6p��c��d��}z3}ǹ�+�f\w�:�(^�t���^&�i�b�c�o1�d���;���"Sj@M�6��A%�j�Gbo�{p��	E�
���Yѻ����	b�pg�m)^��� &���=��ݒ2��i�]iH#çؗ�W�W�h%�0�3�5�]1�M�
�1�dǨjPDae\EW� ��Jn���;X,�c�r5Z�j�Q7((�U�a"��'����*l��r	��Αa�W���'.N[5+�S��xb�gz��&W��y�F�� �:0轋O��8�C��{�u�F󱚶JK�_�t�I��A����<G���[��Ѽo[�xV������5Bwf��`� c�P�@NC�AF�=�}d��[��\^I��@�،ou$򧹽f��ոB���M�	�Mdj�:���	���GRwj�`vq#�<:B?]~qۛ��9���@� I��a	B���nM����6jSm��"���W�GG'1f�RY ���;K3�<�M���~S�����T��Z�O#��#�A���~m�I�A@kS�Vf�Ʉ9gmý��� ��Ŋ�=�V��V��'��6�k��:�ﬁe-2�������f}i���������*�����v�߫V@�p�z@	�c{�J��%��F^r�C�)��I�VJD�y�k謇���M_�5��g��S�y�����jK����*X����P�!���v�m��J�F ���x5w�0�e7�R�=�Z���n���EJ��!�+U��d�'���
��r��F�y���~
L��Vv/�!�֦/��/P�W���$$��+,�]2q{&��5�NwVT\��`�]z�=��5�s%�l,�t�S��
I�'���UUf�9�
��4E7d���?߳��q	>�rE~L��kE��eҸE�h��� d1u����Ϗ�X˓+�e�F�-���G*?�u��|��qग�v�8>�C�:;��)�ص�uvs/no��s��t(P?t�>�_u3,�i/fv�l�̩��4SĲ��Xo3�@����Ss��OC�S��ДX��J�Sa���;���F��d�S�wS:�p��Q�ur��A�J0K��_1�{j��d�;ޛW�W�z	6œ��j�·k�ƹ/T[5]P��F/��ǏSd1YÛ���V�U��\��ʓ�S�u�-�d�����>��.�!��o�e��톶�r�5� ��M�o�+�c��z���M=;��<wGŷ�j`Gr�+��i`E�}9�W��jP�������7��^� ���V�RI��X����bΖ��]<D.chu�oP�	i8����+G3�(TSUE�#yvRc�����:��U%��_ZIϐF�9-
G�X��[^'Ę>�x ��Pʂa3m;��D�+�@���bP�] R�%HuHs�Xs������zb��Q��: ]�
�yT;Je$2�	���:3LE1�)����p[�[�#���(���ڭ�GJ��G=�v^��*Td��˳�*�/��(!� �"�j��x�Q]q�6W�4+_ɀ�?|S�*�}����`4�X6~Κ�g�"�Ue�X�i�U�"tj��<0�?�$�����t�P!�pM��1-Ul̛�� ��g�/��c%��Ӑ�_�F�\C�|@B��9�;"A�c?��*>��Ij��x�X��ڴ`Z\
<5@����L�Q�ơ�uލ�m�W��� Ꟛ|��@(��Ϋ�
�1� �u= �G���[�5g���������(7~� L��b�dE}%�q&��;h8�,lW<���8na4���f��5����[���|'ִ��s�?���̫����c�סޟ�MN���-ۈ`����/���P1M�x�j��8?f�)G�ay�g�x����r�{vZ̞&��+��IO�)�AX�X�גH�\<#H���G���<m��E�s&�wg�T��Ȕ~N+<@H�zA�\��OL�)������[�=uJ�0R���'3�f��*���mX�&&��-�Y��8CA���m��o9X�>��6t~7�B�<�����S�N�
��~ò�������DxC?��QAV�[P��E���F�4<̛3 ��iM,����ۄH*ض�ۿ�t�v���!�0x`q���-���ޱL��|o�q3^���l?"�-_UF�*,��hk�x���g��J�CA��0��I�Z����Y��}>�	;#��4{����{Y�6�G��@�nMЖe����Б�e(��0���0%.�����<))������+��}d