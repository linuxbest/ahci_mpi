XlxV64EB    573e    14b0�ά�4���!m�\3'W�J�h���z�'a� �l>Y�.��`��Q��D��&Q����y.5�W��0�����5S��s��6��"����S_��a�7ݜ�l�S-G��є�$CV1�@k!�멸����(�N�����|%�/�Ǩ���:R����C��Z\�`r��0��΢�>Oc�D�e�V��/4f��;����"
f�ָD5�/Z�C��Ū�������c�-��3��.���s�a~��.؛%��6���ag��{W�PXF�f��끤+���%�&�,�r���xI�\mU�Kґ��n4,�4<�m�74�qڢ��������ɻ~
��6_H"������ѳפcd�$D"/����	-.��?�ڇT��!ՉޕB�Q�>o\X�X�b%~EK�4���nC3��'�')i֤l⑨To�F���k�2C};M;�|&c�q��2wd9���,h�����lp���(�_i<F��5��X�l`��|�I<�Ƃ  r��V�l8?��i�݊�Hg���AT!����Ek���kl稲߰m�|b��M�C�~DJ��K}���� ����qW�%5%(�܅x�KTk!����)l�ip@����%�٤��73
x�UŰ32¤�Z��rx��� 紽��T�o�d>F$�!m=2K9%�����qkvڰŅ���>��)�|���]悖R�.?Kkc5-h��K��X���v�8B�]3�c�����?c7����y�Hԭ���� N�ծ��.������nX�1Cᯗ��ch��JA�q���3��"�ҜVX��3�m�s_�Bє�{.���u�fo/a$k���k3,s�goPz�pVF:�\DLwY4��uQ�7�\��E����@Q�}pe���j�k��U�� N���*����΢���s�B�GPOm ��¤Tkn>��	S�v�v9WI��X��M�ŉ�4�?`���P�8��:Re=J�m���D��m7���T�g�6�u�5IB$��$�W�2S-c�h
i��/��Nm�!�g �Iyۊ\Sk1��䅎�k��CS�?2Q~w�G��gb�9"j#Y�"d!lW(�5fC �&sA���Y{h+1���u�[���s ^�5W{�e|�����qPi��(H�5}�;<P��'�>^3��[�����D�N�s��ى��HT�ʖba%%�X��i�IM��[�)��މ�|AF�tx�s��Jǹ?����A�1$2� �AH0�hv6`��2S�=N%Ҫ�J��-�akX8�V���`��R��v�Ր����O��0�[l2H��A�|���Z�/'��qYW��ļ9�)^�(�[��K�|�`A4�ߎ�����2(���ş��H��w�9c�6�W�����XI*p�`��u���,*�V�t�f=!�0&K7��;�x^��ɦ�C^=���uz��x./��'���*o3���ƘJ=�I�
n����_�7*��%�z'�q3�3�����w��q�4YY��"�i�֦G3+�P�i��R�h��<%���r�/riN|"��[��x��=�L�dξĄ�7��a�ص�~��]��e�n�A����;�EC��h>���-5��)�o�8s	b��pn��F�'��QJػ>:�'��{��HWr��?JM�:YT�Lֿ��C���m||Ycw���y5^i��n�"x#��~~��| �n�]�c7#n��0a�h��hG�M�M�6n{�ҩ9ROí����r����X�&��7:��\�;����<��{Sr����������g4œ�!mr�R%�ʝm���$mN�ޣ�����B�ɖ��S}4�����(�^�)�@%Z�1��y5kZ�6Aqӌ�izv���8�C��ݳ92�j�$nx�q*k@��)��F��+
�^�P��� A��r�^��t(�CVn��S�w�P�F*�oɂ��b��9Hs�2��d��j��S����C�Lb�N׃gB�P��S�[��G�F�zK!&�g�B��t�D2�ٹj|,��T;{d̈�1(��1a�B/b�|�jEħ�l�Pkz�'��)V{��(�O�_�uLЙ��k�ƵE��GX ^���?pN��*�g�Xelȩ�y]ڔ�(h�rd�E�0P&՘[,�i�=
H$�#�?5[���O��'�l��-����m�ν.��aC�{�'rdЀ(���ai	Yt�ZeA����)���!EQ�I/� y�=�p?��M�#��)ػK8���F�Po+@-"��^-��UL�@P��A&�j`�M��K�����&�s-bPl@@�7X��Ϲ�T�H�9a�F�g�!(�����������i]�`%�[2EKd�rtV������c�E̚�$��Ӵ�W�f��A�hJc8Zb!�p�KA��k�
n���q�s�)�]��Q5R���H ��+���aR�qB����gJ�j���C����U�l���#>��B"���,�2�ʦ<���ئ{Ot��s�İ#qg������_o����s�{�&>�k�M���]��H����I�
 �l!�هf�gk4[h�ǟ��l���®�؎��+"�,���N�Vu�ЙaB�K��fm�͖��ܾ4B��n`U���q+�����y��m��I##�t@&Q�ߠ\��6���7U$7�|Jq�MZ�kY�"U=����?A ���!�J��-���(zSjD�?�v'MM~�zY�巀%Uui� ��(o#��(�P.#��i�eʕu���Z5}����T[����]1�{�Nr�u0�{ק��=��Í����֤ӏZ`��q�h*H����c�n���on�vc1�K,����Ղ*fX�
��C��>@&^���ۨ��#�S^f4���!?�>"7z,��Ο���&lNk�: ����"XSdq�>�2lc�^#4aNH�*��j �5�.����#`}3X��(x8!��g\
���Y]ɰ@����sQ��cvvn���m���ˍf�������<dx�P�h��-��x~X*b>�UV��טO�g!�Os9&j��P�۔�~u^+�����# 2�R���UN�x���O�~�h<���i } �?���|Y�qZ��i���A(��X�{�맘{u~�Vkɞ��w>�������նw�?����L2�ë�=I��Ŏ��'{�.�E7K�FK�����m0�ϝ����M��7��8c�/�dc���LY-����/8��Ϙ\qFn�)�)m��]�N_���eq���Jz�,oB�|�a�l������� "8/q�P�9���%���@:�lL����ȉ����~|>w���L;4��URJK�t������#�� [�Kk_e���`�8\dR]�Tf"d�@ۙ^�u�����7�IY����l�x;ȆP�*�莿��۽Aث{�fz��;��5���d��O>^`I�d|!޴H�AY�9��ư�*����ԇo�8�ן�v��/�����k~� �]N/�)�=�����3�?�r,+�HKr�m/�L{�=�L�HH�
��d�*Jq�K+aR�K�����;��Swo�α&���\��	u 5^-��~��Rv��g�Kp,y;�nIϲ|����h� �F=vn�`
�w�e@�����*c���,���G�i0|�R»R	�*�h����C>H��]�Pl%Ur�W��fkQµ�{"�T�<MN�GX �C� ���g [�K��j���;�ȅxx�x��ǭ�VF��|��5��3���Wzo7d.9~��S�E��Xެ�}����$�����
��=���8�����T57w�c��ĺW`�;k+C	)#���w�b��ʱn>�wǧ.�5�q�J��[�����QDɌ�=��{�ɤȞf�(�":����9��j�}�?��xX���	gA+�,=�T��>ʚ�,�=ox�ը4z��]��!H��n��|����³�V_Y�"�x��|$���#C�$�&�U~���nڞML�NT*���w>���Z�h�Tp�a:jtי�������Xo�Te�<	�hy���beC|��(��ƃ!�N�j`H[�;@��S�3m�
��W4|U����f��̉�r]���<�O�n6��Fr� ��Id�h����@�@����r�~�g3
�!$J
Z:Jh��8 	R䔆�QE`���@�ܕ���l�#pFԀ'��U���:�,]+��$ݧ}ļXK�F��J�?;5S��;Qg'��+�(u\�+`�
��rV	�@�]��oG�G���ڽ��I������+@t6��e��p�,j���[j�L^�Y�G]�Q����Oz	g�D�������g����� �P��F/�kO�[08���6�
�LkK��͡C���qm�u6%{��p?�
%"�������RB���SB\D�g�a��<�{[�-¡�Z+z,o��gl{S�dyW:o��OY�����]����X��6K�ؐ���3\8�?C�Mf�S?U�/Oĥ��U�Y�C\�x	o2����>�Qک�#K���3�D�s��}
x�׷D�!�=�����1�)�U�]���2XM���.�
:�w�$�`��Ĉ�[�h��u>w�8�y�Gy���� ]�ܦ����t��o*�
���fu^b��M�s��}Ǵ���e���m��r婩�#l�!��0��2P��2��ਹ,��|�_m�;�6p�H��Q��%$�y�0�����^C�0�.~b���D�K�9���EZp&E[]�e�k�u&/X�e�<�Zş�P#�-�љ�o� �}�Yn���hک����.Sy���X�pn%�m۳��ֳ
^��Jw�)+�ǾU�Q�Ti���Я7��Q�����f��h��oZ ?��Z������kJ�|�Z���X�i�Ź��̑�fk�JP�+[�����W��g߰�\��2����󕘨��������0lhǁ-W
����)�?�j\�&�-i���H�=wo�f����A��R7��z���?v��iJ����?
�w�4e�H�|�U�P3?G��Y��F$�|f1T��ܓ�Փ�V�x��_f���h��O�%B&��@[!B��ͯ��W�c�hhG�(��84�.�ǫ'LQ��k�U��8[E4�Q��Eo���^Mkŭ�|9��Cc(�T)2�|$ؖVA��ae|f��e��VQ��v�\�=L�G�o#M��̓�n�u�<�q5�u�C�u�