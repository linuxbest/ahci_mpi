XlxV64EB    57e2    1350�<��0[�bV*��}X	[lni�p�TH}�>mG���C�G�m��3}P0���GeI����!AS�S��9�}Exղ�Uv�{9A0 ���e�@$�J�I�s���� ]@�i9'%�~|�|44���]3�q��2��t ��[�?3F_�B3�I�nK_QX:��1O�I�X0- %�>/eb9�ց(��r���?���u3���іa�bD�҂�ԣ�����������Cz��a��6��g�dq3.� Չ,�O�D��
�����Gk����?����0)W4`��x��K����L��1O�&��1����_�.@[�}��w���^��u���7�ȿN�LH"�1I�V� 4l�.n�u*�	JN`6��V�;��v����� ���P�ap20�qC�h��w6��m9RcY����%xb�x�/�ÏE� ��/�8�xeڍT.<<4�:ڊ��q������ƣ��wv�ux`�~B��#O����ƨm��Y�t�ˬzy7W�_�a�Vrl}E�uٚ��A��xO���H�t�|k��0�0��,�c@0��ɢ�u]6S���h�ڌ��y����r*�(��-v��κYB+%C��ۃ@I/�g9��K�Ӗ^��,���f��9Z;�~GT�,+��'�]��I4��Q�L�ON�/�^�wK����L�����>���K/3[ԅ���J#���D+Y��u$0��𓠷��_���ݕR���/����h�`%[�MH��|:�Ϸa�Q�����N1�8�>.6�`m�=�^F@y�~+���w��ӟ"Fy�����@��T��]W����=m��6���VW$�e|��+��~�)nb'��&���Z�X�L����	�}� bP�*�u�\������� ����"g����A�����O����MJ�-> a+3�&:�hHcaO��ڛr�.Jy�nP�W�+˾d��W>�=E
���Z�ǥ~��J�7
�=�޹7�;��'��b�Yk��y⍠��%O�^+�X *��˜+��C�}�~%�ʰ�e(H��3�z\{_��j%ҫy2��j�h�b��Y1aՆ-��ͽ2��'@"���3�-1�Mޣ�j��G�ؘy�(�#�ɕ촾�jn�>�*s4_ӵ�ö�[�P�{��� �ఏ�18�=?*�c�	lq87+,����hz�o
��Uf��T��g���o�_BQ39�[
��A�N`n����O�!*t�4犄Е��Ĭx�*��ZoVA$
6�A�Q����(!�w�zh.��_P��.I߁���܄�9J����v�S|.�r*�����8�Lw��MA^n����T!���_�C�ȗK�G�hp{AU����d�O��T��C��RY��r��T�'ŧ�60���[���!w��L8�x��NU��S�&�Fg݉[h���&��V�O��Y`ޣ"A�1'mhб�)�	���hh���*��*��J�4�kb4��ofC݆i���1��9֋*�P R�+o�� �dH i5��M㥶ǚev�.��䈮�h'��$�����VP�)����`�]K��@�y���U���ň�m�~/eU��z�oZ��s?A�ϛ�$9>3���[�W@ߏL�eES|{�.�Pbv���nM�Ȫ�FVd���ԍ���p�K�+�U>Î���#�&�)hoE\R����aӉ-�{ ���K�V���~�������^��l��"����[��n��8Z��d�5��U�t�q�!}��]��n�f1n(|�]��l����YwB1;W�x��]�"Q� (���2�`�3�$t�h9p�}�hvP���a��vB���L��es��(��k�����g���^˦m��QdۭMIVuI����zA���},E�>9�R�k���L����8D�ڸj`�'��3�]O�\k�Π�c��Jl���f2��T�ҵ�R���k�v6c��@M ��Q�Nڟ�a���à�@=�
�b������ͨ�����L��	�=a[��N�y��.ɢ��u⢹˘�ĵ��SeH�ȍyI���!r�n�*܏��p{�e��ȹ��_�����4��8�T��e]k�w?H&�8HWn9qa�2	�����so��k�}G�`!�1���@�6EM	)
���r�0���dږ�N��II��r��#���N��=ӥo���Q��:<t�*.٘s���?��
��)3��{�z�CdU�����6���a��T�n7�k�<���'�x��M ���|cC)ot["�Sk1+�b��MeC��3�њ �ˎ ��ģz�3��F�Ղ
h���"�d>�<�T���_ṋ��0���hh�����Ls9�5���Z�$ʹ�NG_�k��?�M]�8���(���\}I�v��T�G��J��.@������ӢQ��1���z��ς^$na>���o�	���6]�˃\���
��盇O=-F�vR�F�	��e��3	�_�����o��6�gң8X ��>����[���@�&l�����"b��s���d�)Y�hL�O�־�0�>D�L@_�����oxzm�ba(X}���v�1���+���]KJ��37�SU!Q��Dl?z���8a1���c����Dq�i�i`C�?���^p	���78��B���-��5�O@��O�X�;�1G�r���f�ݫr̺]X�mh/?�ާ<�+��� ��Aݼ���VX0��G���W��( ;)1��l��ڹ������L|S���`H��X:?YE"���c����؜:&|9(�QK�,C[�TW��?�1���s��ݩ�Eἶ.��M�Sj�bK�${�����Q~����
���0��c��� 	C���������� }�		C�uz:+u5?{�\iZ<�EbU�P��Ż}^���1&{E�6�q����
�Y;r�C�x� -��(�9��|�p��a�������������<I�;!�2����ւ�LyC�#�VƼGNv�i{���Gl�#}��;��ώC����v�p����]�m8Rz����76�NE�����i��b��c0f�;\��m��Dͨkn�3���ښ��E��� ���,3���:S D���܊�!�R���:ĝ��Н(<jqiI��#�I��R�_��O�$�*"!�������}g����4��yAY�⢳|���ǡ�ǦՉ�i����ܢ߭d�uI�!lP "�4���ÂE�LIg����(�R�1;:<����G~+�w����t�|��V�s{z_��bM�g���Գq[tՄ�d�d�Lę8P4�Yc~��q�YH1[��:�	u���`���d�k���Yۣ��D'#,�W.Ô�� ���"�{�! ��:%�#99g� ~�k&AwA�΁n��(��FT|h˫n��~����T˽��E�;3iL��7z>t��$�87����~2����:H>,\�vh�$s�N��r�����:c(�\���1�c�>� ��e���r��u���}']=Ƶ�Bk�%̇0�b
~/s�ذu�Ȕ���!=	��(9�Z8�]����}�TC�����+���*l����US�8	��hp��߯(�X�?Q�㤱0v��.d�ѨI	�!�k��>@`�x��
p���	�����U�I���_��㈊��@n,G%��j\���HY�`
',��c��H����k���bn{o��j!�ɑ����nr^L�f�B�%��7���cj��ߑ1�f�蝮1 ���-�ܳQ�Ė~������]n�_�p&ҞgU��9�B�&^:�������;�ϳ��U�-��Q �`Q��=-�>MV��n����p	h��N+��Η|����#������xO0].!t�����{>NM�Ї`��B�����8%�|#������yQ#����z�ޚĒ ��sR��K��g]�VB�0uE@��S������L�y&r�uH�U���#[���[ט�MjV
��O5�E��^[��i�T�I��=����>�࡫��a'��b���w�L"�˴>��FUqb�X���Ia�Q��v����(�>�᲋��,f�o'��~|�]Қ���x�Z�=C���1����`�|h�j�F5]�􅣿w�f�O�i��8�n�ρMᝄ���ഠAB;5+!�B�T�M�Q�T
8�Z��[�o�e`�%�C�40�a�4�IଦdE�!���;f��q�Ƌ���j![�^J"[��5���_3�:���7h�����>�y��<���r�VVU�E��x��(�si3����e�U�(�]��A�E����?g-H�޼�&2ƥח1�a�ϖ�"��"m�(�@2U�6�Y;���j��L�@ͽ-�ᇲ�!P�	��y��y
��Y�~��}������K�:T�U��'7$�fd��'��
�Vjb�~E\�k�Y ���Drw0oJ���er�1v6ґ+��eM|L��g��t$�#
����	�y>M���������1m�%t�u����������^;A�z���&�M��8aGڵ��\T#��p���@^b>AK�V�S�X��y�W,����."��h���|;�� ��"���lKW��E7�l�ox	�s-I���P�x�� ~��^%Y���̫_%�@TkժJ���>`�������GG[�r��䓗��{�\_+n�nՖ���XʉY[a�٭ne����@�4�Жp�"�Cc��|�[��
��#�,�E_'u#�!�{T$�E8' <��Y%���>\��/]bG_�O~	�fA�_��C��l�m��GP�/��#c]G7��`W�{� /����ʺi r�����iq�G@OEX-��{