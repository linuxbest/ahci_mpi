XlxV64EB    571b    1300�p�q9�u�gB���<�5���V|���.E�)3
��\���j�201,a	�S��wۈ��r#�nt�ȝm
$!͆�e����יE�T5U{s>5����X!xӆa���C�	�_O�����:2LH���tͭQǺ�;ֹ��������Ew2R�湣!s��- o�c�K�!��M"HQ���{��-��Ӿa�ūM�Z�z��p��7��y�^0�<�{���B���+q��*#>'3!����^��Zl���u !hx5�pWd]�.��F����
`�s�!g5�Ӯ�X�k=B��¯�������;�B�BFZ�ّLq	�?�FL����1�?M޹	��7)T0Ìi��]h<)�2�_�i-�3KP3��D���$3(��aҘ	�.�Ђ]����eH�+��:�ײ�����=5w�N�uJ�ܤ����]�9.Y��j8@I�ӈ�b욷+jn|^a&�h���a�WpC�F�1���z�K������:�:i��s�*~�.�����0�)�D�x�갛� �-�� �=o�/�H*��n�o�4��|�ݶ�E���As �g>�����y��Hs��PAW0S4�Df'���W������P}�oq�	���P�,b�3�]�[t=�^�s;�;2§Â�Y��Um�� �5��{����# ���.��ڳ_|���>1����f(�_XA{���re�Gø�E�/���A�>O�Wh�0È>y�������閷"ChT���/x�����à|_�/�4�C�S�-����W��K�v)D}�g�FH,����!�ZoE�m��}Ẽ0*}aa|��1����BA�����`&��q���繹�qO#�A�;�Dq���>'<<��f5�D��F�>DIyg�#$>��B���]�2��=ҏ�,	���MU2h1:/喞T,���X�[����Ĕ%m��]��$́O����o�W�i���ɏ)��"����n����ש
��.���@�_L3>���Eg��L=*��f����ѹ�}�M��|��F7�T�w_����9fe�r���Qռڧ��k���@-F���;��wȣ��k�`{����ܡ�;��f!�LP�C+�{�r��.�C�[t�m���@^h��|�%�����v�a(k~�����(e ̂4P��-��Q.,�C͉���I����Sx�;Wx��*��a���z�����Ԯģ�*IpG��l=2�^-��&	+^�b�r��3(tb���ψQ����nr����}��*��f&�tX�}�����%��jA衍~�eDk�n�lz�����y]�/?}a��sWYd����7)\���B�.2G<��!��j�:�d(R?��h�Xû_U��D���Y���8Yu*.�2+������Ċ�������t+�B�`�$�Cs؟R��]��Y��V7V�X�r�}Cm\?�g��)���>_/��c����{���u�G�-�ӯ�"Ae�L��]>�5hm+�� ��$�S3�f��ˬ�Y�����H�[P3�2!_�x��y4��5!��i�Э���z��k��7��e���
��w�"	n������W��R�h'\�J\��]	�<�*Y�N�x&Af�9'�%;o_���,P�����tGZyg����p���GR�4�A}�u���*�8��܋�Wc%�n̼�d
)Qo,�+;$��^�wg#@��Ç���Ϥ�ݜ��MeP��%+�
��}�����q6�j/J�{1�]�`r%}9��[�Ā� ����7���O�_�M����ޮ���3� �w���QG
�0)E�-������v'��}b�o�.��t`��t�t��ůé�*�zo<�K�
86{�{����w+b�Q��!��V.s���`�϶Y��418u8ZT�|�#�_}"w��>�|�}~�����h�ș4օ�M�������\��=�^}&Pu��������9��TM�p��S�C��f�6�B��Q��|�Ov&�/�hu����^{����M��5�w���%��W/SE1�p��4��~:RE�r(p�k�A�>֎���Nr�#�i��4��1�(i�f5���'�\���[,ƔO���U"��������Os���T�X�SY�EҮ��Q��������B��4�����J�C;�������a��j��t]�ݯ�rs������k/�_�8j�IMaa;�j�6�?D����p:���\n-XVo
���h�VV�bT5I�L�Tq;G�w	�!���D؜@���I�<�0'�x��M�!W�8J��C�6�}�НM�:�t�{�'�.S<�B�9�d���&m�����(%���M���I����6ر\�Mߙ�geɪ@�y'C~�d�㟷y��~i5j�C}��%��.*h�Y��zU.������Qi�M,V%;�[�V2�UH��|�Y@���)����-Ļh�wj+\�;ά7���f���P�ZO?�2?`�2�[���q�)=�>)1��A���.���@�0�:��n�ќ2�=&�&�||�W1K�V�a��Ѕ���f���fl��x��f#�`�!wa������@��pa+a�]<G[A^�����<� ��9�n��f�T��h2���}� �V8��p�������->k����j��3��r�O�Ŀ��ж�3Wؒ呼������R����n怟�+y8���!�h�RA4ɳ�<�+$���L]eM��x(j:)���T�[d?�+�#�g���EDl�J5p�^�+2b�a�՚!Iu;)ǉ��ټn�Sz7ZJ�a����.׾|��U�&�=czY�<�LS�R'W~ޯ�7a�zxE{)�-~�>��'������r����M_Ƚ�1�7��/��C9+��r��u��WY2.O̱�7ý���� Qݴ6�4j�QN�J�C>%�I��l���[�ͳɃ���d��jYK������q0rZT硱sM
�A�X>��k�xrК�_��h+C�F��\Z����#Dҿ��aM!�z�w:1��)M�!+�=xS��l�ڡ���W�>8p3)$FҊń��_]U�p"tM/T>�T[^T� �E(�$����꺝,�����W1�i�b��7+6��h� p8-9Ca��j�� ����Ռ��w���U�TN��jѝT�T�����~]�ָU�[�>H0s��� G�B�IY�S<0z����b F��P��	����G U!�⯂L�
ivC���X�r{Wگ�;�TJ��΃�;���,�z�xA�+�*�S\�$�=��t�	��z�y�R|��̂Fo���t�z�a��Ki�4x���l�}=4]X������^Նx�^���k˔�� ��@w��s�i���n��@�����D�C��$ߗvܱ ?ɮ�=BT]�[���EΞ~�[6�^�3p �{0o���M���_�Ƕ��72��j�����Dc�j�����A5	�����"A�"�yu����3+�G�Γq��8l��bp�����]��H/HQ���:�_a*��o����>��,GE��N�ic@��J��qg��PZ��ɕu���3�V�H��:�!�
�5�]uDۤ��q�8��؀��dH�I�q4��LGӣ�]�q�5A4��Jx>>�H�qS_�d�8�����Q��1T%l�B�O#>58j�ENи�n�j�\}��
O�!�cg@^�������V=D��?�vQ�]1�2 \SݖFHV�67���)D`6����_������"75��>Bz÷��.���q��[�?0s�����+r��^a2�ls��h� =��7����8�8���w�4�Cʐ��S�
H��jM�������Z�kr��uAx�C
r($>^y	_F&c��|�����6�v�ڇs���Oo|�	�..�C�i�gY��@���+�������ت ���/
���l>*�f���'�z$�OR���Tu�ʙE>��0��$Ϗ�A��e���4r� �ґ*��=����n��1��'_n�u>v�@Ί���R~_8�J�O�:tC���xC|<�A,�A��cɔDѓ|ާc*y�bh*�ks������1����4���z�c��:IwD�|(Fy�d�&M��B٢mM�d���T⻜�j�G��� �~<������U���D6�%3m���)V��Lo_M�B�)����}?5)1�2�/��5Rc<�*b5������-Ψ��#e��{A���̷bd�4����Q�'�r��up���"p	�V��կ���t�u\������Ơ���Ð9�d��	����r��K"R����jT�˖<i���iLe.�L1�7�Va^ ~#�ّ̆��x}4<�	����씻�;���^�[��T���iSӜ�V��P�j�gv�2C�<j�aWZ0��&	�2T�[�K�{�{'z閻�䙁��NҾ��2��L"!RI�v�V�v�ῃ�{���T1:��ɏ�`�M�r�._Z/
���|�S�#M��y4���m6x���G,������<�л՟�+�{3?�I��!��kl w?VI;w�|�p�	7'���63њνŴ�NM����2�N�C�1��9�� hjQ�B�K�;�0���%A�
��~�L���z�/���n���A+�=_���!���Pn�Ϩ�@���d�7Ȏd���C��$$�qh{M��C��xXk�U����{��|��&�:(��_"��}����$��\�F��& ���EE�J��V�Av�SB�< |��VY��ie:Ȱ h�`��0��T�k$�6�ּ	�1p: