XlxV64EB    fa00    2c40P]m��
¿�O1w��T
5{�C`�=q����G���������xy!�����pP��J�v�q.Zwy ���1��X,�Ij�\$�v4����ඕ;w�XLX��f|3�>���N��'d���=�?�25.�&m����Πr,|�9#�{p��o|�7&�&�\94Eq��q	��i��x�4�ۓ�v��H�T[�p�6�Y���\����s6��2���o�T{�CԚO#���p�J��T_lӽ��M�8�"�'z��D#F�^@�P߅���sV�_h�@ ��0V3D�!�88���N��8��s@��� �2��Xg�W�����l[ �HU��EaWz[+�N%�8'��4��TV6o��B���ؒ��#��d7V�$�S�xK�sE��AV�� Bc�d���i�}�?�n���E�[[2�߯B�@���� +�a�	$ԋ���G�v(R^l�ney@�����ߪp�#qH��)pI�� $5	���!��h�ߟ���\i���r�*���}g$6��=8�Yt}簼�$x�U��XA^��P�3��tTR!H��u�eN���B���3�2y���PΆ��������l���V��ώ�J���6�'*�6��,��w}{���R�ġ��*��%�9�s)���'��ł`����ړYL�/MG���!=�_5byY�c�w�N}E�?��8�X��	��nh+Tg��]9q�9���2}l:&	���8�?���aEb�$�4���#���#�Z�'��������]
8�tA=K���I:�v���zB�ƹ��׻�Z6��6w�2�ƚ������nS<�������MT{�j�j�9s��:w�L��T�x���v��$�.CiF�A�I�y7�-8�L!m��+��W�b��)�VF���r�T�c��|�[���)ˀ�������*��?�Nu�b=��f�#V�����鶪�*�ƭPϖ�o���	�*qY��s� #t� �q(�1ӟ��^����0,���!A�j��||n_2��ԍ��/��3v �$�g`���y	�7��M����U"P�oq�n��M<��IdsP6C?4�l�����ݨ���ڛ�3	H�{{7I@�	<��O1�s:�Ű��v6�P׸
SC��}Hڷ����}�y�l
�g�Y�a�WXAk�M0���0��G����^��
�.pSe���8��������)�Q0Գ����+�u��-q�m�rP����瑭(M2���M6m�X�a�CJF��u��X稺�w�(R��lu��^0��r�w�-��r�]i�%ν?���^���{�A�+ F�{���5Y�F�GE�{"�@;{*\X�5���ͻ�SCЃ" ���������א�T)��֦_���f!n�E9ب�>{V�9��N�c�<ѕ�$o3��w���X�(�.�p�=M4�v�!��|Ks�N+a"�&?��Ϟ���?��Bv��H?T��TS��v�w@e�u�/�Eq�7��j��c>Q�~yҤ_�c[���;���5iZ���'{�>���!�!|��̗�]��RFg�_����?p�C��e4�9C���z��`��fDD�VB�ғ_LRsGo,��uݢ0���1�ĉ�nU�7L���;zZ�D�Ȱ��Q&$�
~Cl6M\������T��_�I��E�uQ\�`�ْ�ނdMY����;�?t��K #S�9�����L�M"��n���O��V�`��:9�dQ�N��}�T�tٚ,V�&�{�t�Lh�.�PM;_qj��C���:�4]1�����c��"J7�����V
z�g��	;ۅƧSVg���
&櫗|������yTX��`�"�5x��U�0���v��2�eI��Zp�����u���ZI~#=�(P��x�����j|�"��7jօ� ^�QL�o�_ՔU�ND�\�`����.<�d8�5c(�o�D�����pB��.UɍDe5EeHr�NuH4<�+�|���Z�ÛuM�6��A��$��I���ֈY$��17��ܐ�O���	؄�'0R��/�a�Q��Y�c>89!fX�ý�KgF͋UU�qk&W�+����_�����0c/�+O���G]Q��WRG���B��R|�Sy�ͱ>�7��Hk��^7�O�R���[;��	q���я*��F@V��zn��a=޴H�Č^����v���4��`�#��\����r��yk�j9%f��Y^�BG2�NAl^1c	�/��9jq����
E�O��Z�Ch��\�"���9뢡��v� 8���ͺf�v-0���$� Wu[��+�kQ�c�q+����$䓨zukB���K��_S��y`��TW�}�Z�I(�ڇ����,���b>^��L�h-�
J!���W�ތ�Z����Mq�R�bl�A�Ƚ����k&���I���Ϫ��Ƌ(6g`8lC�����PX�r}��4X�,����r<� ��Gv9�}�����ԭ�y�;-Q~ؓ��b>b���\�P�Ӯ�ߓ�˩�������	�z�8G���_�������l��#�����[_�Kz](��C��n��yi[���f99a<���a������	Rm��&��-=��l�MU�&�}}�|�K��bD7�8X�K����T߼<
��"ˀ��E+��㵣}Vf�Q��~{ҹ�B&���C�W��d�?���Ct'2+���Sb+F�Ep����xI8�9���%J��^f�
����Wj���Ѹ<j[͔^*��PA��NФ
�_e�>b:��L._4Ec|p�e#+�OZCZ3�m�eP�;l�o^�KZMW���]�A���l`��M�P�'������o��PzP���u �ڂ+I��A�L���c��>w�s��cM��9c�sߕ}�s���X��u��mR�#�-��y�0��i�>_�N��I^I�{�:�Nf���H�N�m�B����(7xj���mR�,	�Q+�ED��Ov��e�;@���K�>���&?���[�m��nO����ن�Mk�@�t�\];�a�J�}�o�p'kZ�8If���.͹�h����疕�i�bxd�z=r��U��s�����j�O@j@hO��T���RJ1Kc!DA3��'��i�����Ž��<{�X��z� ��	��(��5k&���1�1�6���F���7��3�oyr��k��O��L�Dvɫ����I��[�ϱ%پ���e�f��r`����W�\N��B�ԝ��(�.ȍ�e �>F��I"�w�po���$o$����J\��3I�u1����� y�+��.��$4�$ڍ���z�j2W*�@�@��0r�m�b+��"�q"���E�0��D�0z~ L�^�?�ξF��]���.��@ǻ����՗��]�}\�ރ��!�7k��=�^Qq(�qU��j�t`���(�d��
��%�r��g9}Σ�P�(�7�B$p~�/��8����c�d~}@�F(����䈊��h�������%>3#�f!�[�����6q���H�=rb��)�����,��]!��Mf���.K�x��h�����n,$>}�����tg���,���p�	���E �6�\=+>ϲ�&�}݀m�'A=��bS�>��$@BO�5r�ٶ��Ҍ꣡�-�D3�E�3J^�h��
&k��m{q��e�LJm�������!dLGX�j�l 7z�e�X	%us�/ɐ`py��H�t<��q��P1� �e�ն��j�hKҶ�,C���P�����+��!N�;I;\�A�.��XjD�@>,���x�#@�:<��������d������RRI��I�N@��Q#|K��BP�>Xh>��� ܠ�#� M
�,Y'��y㊽��7q��.����;cC�7�oN��_&��'inIug��/�񳪡%�R�-�+�/ ��7[���b$!4�Y�2r��h�Wi݋�+����r�aّ\O{Z�Y�䷣�5��G��M�z�N��&�gS�����|�W�0zP�v�0aC�6����.���9�Ձ����7UZH�U�Ty����V ��ۓ�z4@L=Z�m��:�(F�u=S�
]�H?Pc,Qi�/�a�_�Nf�n��E��=D�f�����T���v�֠�_�Ty�ӑ���ͲM�X�����n�ye��3w����(�+���M�t�T���o�����֍�� PX��M�1��LB����yQ�\(������f�BS��X��i��� ����X֣M���c�3��^�!J��y��1KWu?R$o3�ɘ(�3~e���4��H_ǉ���ˌ7̭��j��hO�/���΋e��p����}"�w������$�K�J��g�F��"�B�N��;�����5���	�)����`���JP7DJ��K��	�.ıe�I�/�-�08�$'N��l1�j �4Х-yt�ܤ�N�~�Spl�󢌶e�?_@�1�˧Ɋ��n�nP�'�2.g�p{mw�m	�9J@�G�,b�n�?���y:6X�$�
ٮ@��M���gن��!���.y��Pw�y�eeM�'�3�g��n
X$J~')9ڳ�F$�QM@�t�@���E$�*��}$18P�wY	m��&ғ*�4�<\S��^�;Z[�?À�M�;�d�#�|-��A�����?���H��Ԥ	RpR�-H����t�m�P�]_8���g�1;�!B��7���QJ߆A�o(�=��/��FL�&��a�RB��t��3Z��F��u��������a^x�Q�`h���	�a��Lj尃�V>k����ҡ�wQ�ҟX�Ǹ�E�iķ���4�۟ �78Y��R���qo� �����{w5m�ξ^��{#��4<%p�{��)����LĀ�>��|�d�,�����MN�؂�@s���*�c�8|�I���Ȭ�'����,�'&����s�
�>F�VA��]��n��āo���M,D_̹┒iQ�M��j�gw�����&}<��6��RӐ"w�-v�#���{B�K��R�l����x�:)f��XzCB�
{�/�&;�C���d $>�4�t��;S
�1��ϱ4
r����8(�~�Z�Z� $����h���L��5g�Ջ�p�wnz��U�a�Dֺ)���p:x���u�0�]͒%qBg�0/��yjL�����$��3y���?78�h�it��#GJ�"�P���"4ꦥh��w�Ņd��U��#�ܞ1��o�V��D��F��F�}�?{����j6��'�!_�7���B��c�s�ܐ:Ѥt���3��ooA�4��B����*B֚�9)Ѽ�@"	+$��\�_��YM\�|�d����=���9�	R�ޅpI�v��	��x��D�qÏ�V
����#�� F��LNh!֢��H���
ϑ���=���k�c�"ݗ�����C�jM$�IP-��?�u��nעΕ�/��D���+aQ� �ϙ@���:�o�Q����O��i<�."�`���x� �?T���J1Ls����)UI�z2����/�bK������/{:�N�I��@�<1��+�Q���O<Y�ED2� E��D���aoMy,~��}�	�I����Er���y�u54\W�[�؁�߹����諤i�u�Sd2�t�Pu����t�}k�g�T���Q�q;�=��9nySf�T�&	&�w�$���LB�:ݭ�M���4Z��&�r,p�������9��,IA��H�ڛ3_?<E��`�x�%':w�;���#�"�}��,���JF�YJ�E�;��ך� }T�1v��[���^FB
[S��Z�� 7nS!e��`6.�_���>������7�|�s8��u����/r�Vs� �����SSxjB%�/����`;�k�è}^L�
�p@�=g�Y���7�k�ÚvAE&��sy�rd����Xib�0��;el�u'iP_��1 ��C�����J�g@V妆0�b��|�DLެ��D�a���5�)ϭˣ��]�m��[�����1p-��E���٪��P�>a E�) �wL��O'>�"+�e�)1.�A�6d�40F��I�5��un��f)�p@#;��b ԷK0OrX�W�����D�M'j�ø��[���An�~�y�@���F�]+�Fd�/���cI}^l�_����eK�#J�\;�Ҝ�c�xU)�����2uB���u}�`y���q��U��g�M8�׎�q�dV�`�X^��d�D ����k�8���n$;%�TP
�e����xDۊ9;R�e��"�t�Zue��}D"qQg�;� �������!������>�%io��Y-�DE�-޺zL�1_c��2�v�!�y[U���"��K99�i�`�-�Y'��� {*�P�	�ޮx�_{O]���[����$��X!��W�2�B7=�%cg����C�R9F�d|�����F;��x�u��7�ZNBq����*��ZF�I���ŝ�~=nMMx��À����)J�>��1�� op}���n��$�Zk�1<:�C��31���=�xV��������]:�]��bz-a��4G�ZEj�m�pN�P|�gq���4Q����D�E��W��r�	*9���cy�?f��C� �p�b"��˛�H��#�0b�x�Q�]�:���7�C]���DpKA�Q��yld� N=}����]��,Uׄc�����dƶ�
��\�@V6��vy>P�����^"Ѫ����J=!-��X�ʾQI8��(P�2��m"��P�]=W�B	?�z�a,dU��	꒒�΀{xRk��;a㸋JYSjh��=���v�g3�k����ɑ�Q��A9����>�ψ_wz��i���O��f�b��A�ajSm��`�zR��"?�z�LC\EE�G������iL��W�/ ���z|�����<\yw	���:Ta$m<L�ͻԶ��Jm}WvM��"���抢�$�3v�wn��-�iB�tDm5$_tZ���Y�����s㘰Ƹc�c���#�A�X!��D��U�V�
�����{/��Aa5g,�%���=�� Drb���W�%Swm����:E���*-�|@<�X�-#�O�U9㜄���.u�|x�k�ħI�Sy��rZb�q^g���[��ƣ��1��B��*���8�ݽ��<[P,�p���af�j�m
!J}�!�JY6��ŨQ����b�X�Sh��0�fhB\*�r���]w.N�%@:&��k�'�<ݧ���t�u�L����+pt*�6��á[+6�+!��5*��n3-g��\(?��VsM,���G�I�ad5����5fC/������<�L��	����t�7ovWi3�ci:��,��/�E������Jr̪�3U�z�k�ӛs��;�s ��P�=u��rGY�o�a���	��L0rz�h�d��u���mPfeіީ�t	C�H���zWCD�)��c�K�Dt�Fc�$�jTޙVSa�F�+Q���R{A��:�hF������*�p�L������S.��14uJKot�'�T���qi_�Φ�ê�F��9)FJ!�Ҟ��빔G�o�[&y���T�A^n�+�a1ghq�֢�$����|�>�C�>Pv��U�.JcN�+�!,6/�i�c�V���B�$z����S�lϵf�$6~��-W}����ι���8'�ƃ,�Q�gj"�Q��ee�RaQ�_
����yx�B���T��K��,&t=�b7uE��Fm�8��*�n�xe��GP���/�}R��U���'p�Eu�E��R<���]�Z	�/�^_ۓ��*�g���NA*N�W�^w��;tR��Ko�*Ј��ڭ}�iJy#�*D�qRi���p��Է��YC�i���C���
�SNҘo�pM �B���U�	�%!�E�� 
�?%��$(�G�����SV�j<$	u� ��;������2���0⻵"���A�$�L�Ο����P(E�n��`OH�M��!X{�~I�+p7">a�5S�A�CL�=��f��V��\VDt�z��.��sH�:~G�X��s �KX�Lsih��mZw�g�^F��+tEX-��m�e��{P9%HUr�9`�m*���Z�1}.xą��ſ��Fa�vj�C�����F��=��R2�9�T�����ğ���da��$�dp�;��U>?�1y4��EWr�a�WY�3�"7�&� ����w��{���5�"�-r�#\ʧx6���4V�g��=a����L�s�=d�v����D�vp!��<���~�F6�9[r堩����֝��ïφ0�I�����T��~�	��R����L�4l�Çz�3��9H����Up|&{5c'�|B"����լSCA�~@	R�1ǩ�C��+9�����u�n��Tx 64��PⶮY58/d����9��<��0��G*c�E�9��lH�h�`:C���j�b�S1��u�e::�<�����7�
��_��'�,=l0៰+��}`�*�m���l��fz���b���0� ��&�(�p�#��6�"׬�]K t)=��D��h����|����Y��"����%�ߎ��~YGn3V�`��w�gI������R?���)�-��,�:	����w�|�����=}�9�qyCg��,ۇ�rB����7���X�� ����l$4�>��<'�P������`R
���%`���hYN�$�8d�7���4߉��ӵ��S�'���3t+�G�kS�2H�T����yZ}3�C�Z�X3�s:O���Rt��O4	���#bH�N1p�B9�K���@�;fÜ��2�W�����T}26�M�YC���QlJ�k���E���
it{�-��}�Y#����@��D�E��i<h�@�Q�7��U+j]�U��FG�2�8�A)H�����l��Ń��o��Y�짰Y�0ə�\v���������}��I𦜚 �WI+$�)2Hi:ӊ�u2k��tѭ�������b����?�z1A2����D����ߡ��H�m	1k�~H�L��$*Φ���p�����`��Ȟ��}l�����S��u���B��߽�3|-~�����	WI���Т��}#Z��Lq�u�`��ݜǟ�Oa�t����DV�#TM��a�e	����!�����E�Q�w��N�1q&����c��{ͷ�������˹h�B��}�>�nT�~�7�s�J�$��p�J�al�v�:�s�y��=Ւ��=�?�Oi�L�]3�Rd&�4��������+�(!R�����q-��*�I2N�^(�g�KѪ|���ړZ��� �8}E�=b�,C��H�]�t�\aNv$_O�$޻Cfl���5�X��½@�9Ji���P�E���F���fjz�`ʧ���7�V�n���+	��{��(�������|��Z�,G�2d�-�Eb8"�9+��.�lo��S�M$��KZ� F������@}V*Z���#�[��T��[�?|0�zZ�-I���TE������wtG�[*�n�6#�����Y1���?�E:�D�kn��}�#RK8���=Pq����c6
�y��ev47��0����vM���T�ӯ�ET��p��? *h�
ؐ+\e���K.i$�f�c�tt��XSϠw�$H �y�*,6��������m?�֊��Z��jQ��Z6=��W�r�Z�]�%����}�7���7!��?\�)i2��t��9+����V�p嶎�ۭ#����,�l�w)ex�8��)�h��?�t���ܩ��,e�*�Xnd*	A!���A�b_n�]KO�Q��:Zir�W.&Ň`(�E�7Q��[`�j�b������]����o�g��A�͏?��:���!�c}�1@�4�O�K�p�G �d��Η�����ՙ�A$�7[az�¾�}�  �nk����#�)�cY
����9��*3�8�X�B���(�[��럣X�F��N�>�p�%���ea��k���%�����r���ܝ_�7dx8��	|+�S�5R�A�P��n���Ɉ����d��d]:��&��[��}�ϠaA`�)o�tC@4U�mhS}��dt>�q��I��T�Qq1�H�;���W��{U2��H�}U^û�@p�\���cV��4]��7�7��u��:'��1�ɵ���ƽ7�~��LSO�D؏�J���B��b���Z�]��Ģ��/R������N�� D^rtN�����nɶ�	E����IY�]�{��m�`,��Q	 ��o�V1�	�b�f�%�B��8c�C�P���B���$��}�5.��;��~w1��c	��$m��Oh(�9Ӏ����a�G�g��k�58Yٛ�_ZҶ���*Y���~c��
`d#���=Id�N��i�u�C1iz�/?\
 8lb�Ԍ���wPΜۖ� N��{ {�A�2��Z	<�� :P$d���,cP��f�VX����$ңK�H��4R��A<��ܢE��l�e�.���{�C�mG�&�@~*f���^ �@`����V�}l�7"R���,��U�*7�V�_��ִe�����v�D�$���F���.�M]�Z-I����S��y��~\���*Pc4'� n~���d��"Xvq�!!���$��x����y���0p�#7�kŹ	��I�o*�A��}<3�킡;�a��Gh
�6)8�=���)ov�hK/�3�t�&�0�f�-ھ��r�[���f�J$���Z��@y���"su�o���U� C���R��{c$��v�I���J��D^���o����䞖�667�E��8�]��G�Wr��԰�µ����<���P��.v�����	EAׄ�{ѳ}�~@�ł�O���H�&UO�e?ŤS�>��ƹ+���=�A�����5H�G9�#�'���ͫGCz�����og�Y|�䦬�>貫�	�*���)�Q�ϫ_P��4<[�rA�|�Ղ8IwOO�[]rqI�4�c�e��m1���V���1T���ߟ�>-,�#XƬ���B�rI/�jluN���Jz��e���XlxV64EB    167e     570���,~���1�@��W�<O�s�P�H��W����� ������D��t�_ѡ�{�z9$`�q��gm=j��?��� *�;�����}ɰx�b�H/H�H�H���ǈW�m�'I��u3��T&��=B鱢�'O�:�WaO9�Pd6�e��[˻t5F}%����6���@��KB�V�g��ç���X�h�-�s����L|�Z�v+)�V.~(�[Z�=��WD��3K��u���J�ĥ�a����Z�%x��t�����h�2�����B_h�3���h�<�gk��-06N��z��k)����������u�b ﵆�I�UX�Z��F�c	�m'���ȐgN��=v���:�_Ǝ^#�[��(6dt,'�#޷�,F�r���~�q�׶�4?L�x\���j��Nl���D�,;��Yd�A��I[��O9�8��C�K0�|h/te�Y���݊��!���������7\�+�n��1Z���	=:suf�8&G�t�AL�ɋ�f�v���H��j*a�Uk�MR�5����̄S࿯=i`��֢p���&�ؘn`��Zg$��W_d�L;�,%6�x�G8l�-&�zX٭Ψ쏕6}�V?�ċ�G�I�S����6[����LO��<#�yZ߉��i���f��K�M�i�c@�a��G�����근x�1�!q�El�����MKM�rmS�+��Z���ts:�Y�Eg�Ե��v�n���ygp�Ol�4�u˫[�2�xM�K���T�UD�5j�-$`�Z��r�����9�ل1�Ŗsj2<���+Z��,��_�QHK\Ŏ!ѩg�Io3����?�p�­ӭ���P)���^Q���\�1��4M����޽н���m�^ݱ��^̙�T3�l�cNѴ�K3�k�/�G���Ldo�adZ�؟q�WM���ХMT\�h��l}*�a�#9-����1�2e���đ��dÈ*}�ۼ�������ś�c���Ϗ�Qb�|s
�>'�j�P�l/��T�J �2J֣�I������ţ�L�C��`��}�Z�T�r2iv]�o��&��Yl�Hn�0+f���م�<��'�J4�UiK����[,Xg8������bQ�H�4��"#d�s?s1�*y�6p�h�-�!W:����0�@K�UU�H����/`Pݪ��f��F��uEWA����m$�J(��N�)a˞،�C
o?��.��~OM	�b������&`X�V��rF�>�����}F�>��=���!(n�B��n�8]�0�n�Ax������ .�I%f�(y{�'�ќ������Z7 ����G�]�����tx#�|��
5O�K��Q�Ӈb!�������Ru�뜛�D�X1�Z���W��O$����r