XlxV64EB    2d5d     a80����Aݿ���ڧ`��l_�un��e�����5��z�/�7�JV�4���H��欪i\�6s^���E��c���� ۄ��g���ᖾH )�/�hY���rSKY�k矕\��bѬQ.4q��(:�Ȱe��e �f��|^��&3�DbdK�;s�+�g�K���L;���n��,��|^���%ASP-�:6}�d�	�ϻ���FBfv�M�z$��e~�7��*K�����V}*��!�Ut����շ��Ly"�}����Siߢ�%���Ik�,�![A�J�3+���p���e=|�z����BgݠG�z�rN�]��]����!y	��y���fԁr��ߜ���*f<��-Č��KJ6��ޒU�N��YG�Y{�v�Qx��I=�o��Be/�0r6!יM�]oJ� �,vG�s���OC���`��c?1 ��4~x�u�q좰�}������b��v����o7Ș���Ix�>��g�-�`�biI����I�HP�5I�)lq�C2�d����?�%!-��J�y5l�M&��l�)�qƏ��(�C���zv�r����Ɗ��D�E]�Y9/vZW&��>�ai=J!h�7���3�!�]޻����.�� L&�����Gw�7�Ԝ�\��|\t훂7�����7�.w���
�{� ��@9Ƴ�O&4�,��������*�G�GlD�1HD	��'��~7�����Ď�({������z�Jt'<���gSC>�}o�����,�"��.u]�y���l������5�,�~����g��!�#�x�@9��8�bJ��l�H<�R���p��M)��Nd���(���
"/�ԖYw�✃��1�	EW`ԹB*�*�Bvތ��#����2�I�2-Z4���ӧ��7��[п�9��}���k��1��@����iש��Ү����+�z���L�wF�b�{4=����w���Dث�f�9:�����H�����C�z�lJN���<o�!��:Y�򚗫���L���������	��~��%`=N�"8��.��n��ⴟ��ϧZO����[I��+������J���'3kI���z´��\-;�GT^����u�?��)��b1��� t�ʒ$�Dy�H�&#�Π�� �eV|��>�B�S���۸���"R��{Z�	Ͷ�jyY��%66lYȆS�E�����f@d�6���X�i�J�O�/�S��_Mqv�BAW{���1�jݭ��M��՛�.�~��7��j����8�����MX�8��R��9�	�ɯ�a���ܚ�:7��GվY�` �k�̺�cV��@��|\L��~F��d�,��B�>Q4d8%�=�Q�"���������j����u�䞪�E�����V�b;��o�hH�èŅ����v��h;����8g)�S�>\�Fl��X�;�~*�1�Bt]�O�Y��8�`W�Tn�&z�@�#5?������KRt*[R�6d5��ǫ����eL�dM���G<�IQ����[V.�>�璳�\��茿�����P%����~]w��rMlJzڐ!��>�Z�v-�e�/�� U���3�s�= "����)��d\��-ַ�Q�<D�����gt�?΂΀�# tL�u��9Y=�Rg%����َ��ڴ~3S-|T�\��I|�~�8o����	࿇V"���eӗ4��녅N5����Y���<|���í�R���Q����	lXT0q�
�*������жv#��ʽ�H�����(�i�v<'�	�˥u���vw�͟� �ˑ%�-r�:p,��0#�Qa���#��ɴͩ�7o���A�CV4jl 1��~5Z��p���p�>����ύ�tt��MԚZ-,����+6>������,[��s�����ɓ��%�2��ߌ�(s���!I��tD���Tc�m�j����qB�%I���q��!'��L�+��R�a��KǗ�ɋ�;�h�!�x{gU���x�\�B�iG|��)o���C|f��)����t�W՟��I�EI�a�pRkϊx��O���gmz<��(�-�1?b9J�B!���ƭ8r���_L��8ƛv�;�{KߠV ���,c�ʭTb�|A8�f�x5K��"�K<ߥ?}BT���%F�n̑��KtLc�R-��NN�Un�~qQف|[��O�;i�'�kB!�h�Xc<��:M���D�_�	���nO� G-^�Y�ı:~��Gq�[xd��JR�m
�����+�ް�+�}BN�Z�S7�*o�R!�W�H��ȘNj��ˬ/:ip��V;`B����5��n�)�?\,5'<�Q6N�0W1�?���4�t�~��H"�4 !)�k�iEɧ��LR��"9j�r���O?�6�<眫�Zx~œ.+�o�PM��ڪ�rDݹ�=G��!خ�O<�V�o�I��û�w$�!x��7Hh�Fd�'C]u�Zz#5��v���mL]t~��������F��;v��I�q��-��iBw�G�KA�៦�)�#Z`�YQ��;�@ܲ�gG(D�_
@�H?8��QE�����}�l/5��}��#�H��>,�r�ӳ~��}�8`xsf�`V!iʕ���4�)�A�`ֻr��$��J�K��� ^J�܀�������2g�b��v�