XlxV64EB    4cec    14a0��7IWt���X%yy�W{��O���%5fޘ'y�KȦ��:`�ٵ$�&�b*+��'��u*2pDy}��b���3 �"j���p&BR�5�[8�gX7@@�G-�;y7�o&g>/
π�ת�Dʓ�S�E��XJ䭾{D��]>�?J��^��B�\�!��#���Z�A���콟����[*���X{���M�����>(&�~8��D|s�R�)�=�?�j¥���8��l�@a��^��å��R�l�BaC�! �m����z��Y�w�Mww(I
�zn�C�:�!SS�1�l�G]��s>���Qq�EXs,�D�Y���`�zz�$�/Z5��r�r2��|F���{1ͬ�$����	��Ͳ����%�"_�Tw���̞�;ٽ�-�r�/ל<]a��&2��$��n
�x����ץ�2����b�
���R>���kŒ��X@eޡU�9�Ur��2Ŭ�̪Թ�a	���m&�\���Z�6r~�i ;�_� |�W �����ZnR�3�aóR�� �u�F�I:>���û^�<�ڶ,�׮v~Z��]:�M/B�w���mqzq@t�EE�u�GW/&��$A~�Gy���T��8�����՛��V�'�L�?����֟�'p|a�+��8���:�;.k ��z0�p E�	G[.��]�>���B��E��M�9��P�Lx	�^�a7����D��P�̬j� ���G�Mk}����+q`�0���0�>;f��25�gu<��0]����0��f/�(^�aC<�"I����{������>�핿Fb�S��c�����ɲ�K���(M�?���fP�s���Ā
�Ͼ�����3`��49u(��nز�Uiz1?Ǩ8��t6 )��C�u��,�����X���m͵�˳8FI������	�S>YD����vJ��$�~Y3'W4��6�5*�Vt���-z�#_�G��5� �a f�ܽ���IQ�Z̃H�2�ܰ	v!O�~A�*���ū�����r�W�d_�r
��vd�ГY�*��~i�	�a�bT=��?c:��@D��_+�oG�@\�	c�-r9^&f�Z�)灗r;�Ta�FsXe�����#'�z��~���u@��x�����%(zΥ$���O62\S}PK��u�t堶�II�WpIh.ů���ʔ�;=�#��H'���Q�,����٫��z���&����>	ܪ̸�C�� ���-�a*b�nJ�}7�sS�^�*��2Y���cçΙ!���+����_#�*&h#mF���s)�U���I�G� ���4O������Xe�T�#$����
�nN��5g��+��U���t�4��0l>zbI_ȗ+xد�����Qt�M*��q�t��>���㙓+9��n�j�^����-J�l�kq�0�q��XD�S�$���"���Rκ�e�뒶I8ڏ>�}�Q�v��AW�*ޕ	֛57L`�$�y�J��k������A�p"�8�@<��b^�w�]�\wvHP0�]��Y���3ū�1x;Ǖ�A$�߶��Kf�,�L��IX�{m<��Z/+�V�+B4Ԉ�]�Q *۠dɊ�|������l�ΥF��b	����l.g����Y�[̐�GpK>ٮ�����	���x��A7�o1Վ�]��S�<�Q�}�����	��A���y�G��؋����YS_��j?�9��W�����6UVU�w�`���J�/>��Śj5
8a��
2�&� �^'�����(���p��y�x������3�G�A��(��C� ��2���c��T�4�,�GkS	�Y
��+��� R��J|�_�i����]�x�d�QU�9�����(.t%`�������`ř�!-���o�x���v�;[�J��1�ޤ���(JWޤ��H�"���H}���	l�i+��}oF���X'�+gC���=�Ϡq{L�Ͻ��d&[�T��O��*;�m5�DK����䴟�}ϗʬڢ�/��7�`�ֳ�I�����L�':���j�a����J�O����{�Q�t��4K�s��r�Ǿ �B����'pz�
-*�5�k��t!���7�ң�jz���CV��+{T��QŊ�؛��i�u1#�;%���pƊ�02L�vf���a[)��ro�t��� ����-fa�mp�uB�4�.{�����z�u����ҹ?�p0��>ܳ1K�Df�@jTuL�bNO���!�$��LD�<"JL����Y��f76�n[�@�xv�cc����I��7����ߦž�?�9/��L�:e�=������k�:��ӈ��R�ܮ������`j��\,��жĆ9"�㴚B���s��v��!h���X�"��$D�X����>�[�~Q�3�5f���pI���D#�2ٰH�['��#�U]7����iHI�LP7��I�� �oZ�
��[�O0Nә��S��1����>���7�[g4�&4�n������Je�r1y�&K�)qx"'�ݐ�'CA_��XX��kj�+P�dz2]��ۈ[T�F��A����9F�ĢV�A��@�d�����lyF���ʑ��<� ����W�,����n��r��K��H�os�<y̖�Q�xzUd��@}��y36BRb�<?l�gJ�����5ZB<5���b�!�Y/�F�zf�UR�:��"�y� o��8��Kr�Jhʐ�}�_�Yhq�I�'�-,�F�������0��*�z���Ч��r�����[����͚�PH��#eo��U��H&'X33�`�E�y�cF�'8��<φkX�*���z��TPJ �5����C2������,sޯt>��]P9��~r��p�'�em�X�:�`���Af"#��"c8?pf2���6�o.��9�ϮS�&!��+���&��7��\��a����$}OamO\��N���j�K�	@:���͵#rd�e�ڇH܆��q�Q���i���I"9��҆	Z��VG�53�f��R��g�Tc�J��ŎO	��_���O'������*Q�=�2��gFi�����1���3�����jh��A,�{�|*}=�\=,�)�J���-��*Na��B���H4 A哩$k�jc�����*f.WN�gXFCba��Y�Ι��3�����Ht�!��:�vp�о�l�l;�|������*U�w�sV]��jT'p�/��ݔJ{�q���rM�m��<(l����3�����K~J�����
����&|�x��E�	A�);�'Te�)�Y�����#������+����Do�Rޗ�g�(���y�g���MnNǲ9|��Һ��@ ���?��� �6ܦש���ߏ�953&�m������[�9�~S�9��h���LU3P�w^;��fo��ԸsK�IX�޽���*)j��C߆e�Ls�# /�_���8�l\�#�����P�,�q�H�ӎ�V�^{�K]�X�Q��w2�Ӭ�7�Z@n���gt��[��bRwG��|�O�̮~��EW��/���"�ofF�,Nsso�BuM���Q`��F�@AB������iJ���3��q��/Hs����@1Z��	�[��f�z�: �@y�[9	5�R�ev<�]��Īц�7rp�hN�궙A��M*�wq��i�V�(G>';� �̃�t��e�ɳ���i��=!%T���������2�+����m8b�unؕ�fg�Ɩ�%~�r]���d:�q��v#���D(q3/���	ؓ��yw�#S����y]���Z7+H��kA?��˗ڼ�,\��*�Ȭ���B:킌�8����.%�9�'rF�+�{h-�=�e�g78��Jj��D��K�C���!�!ms�tG��=�}�D��"����vY롰w��id����3v�c���J���`Ȍ�3�G��k��՚�<2T:Px���?,_�v�G�,�Jm#J�U��?�� Eɿͫ=Cj��

��PH|r8�R�@Rb��I�Ƣ�uoP���uQ*h�ip�C�!�� ��J�<s��\F�E];��;]P ,k8���(����qkRkR�AS�OW�&$6XI��ܻ��d������L����ߔ��Ȋ��sDs�|m�㊩�%Z,8s��EӒ��B���ڋ��3!�v�^b���޿�!� t�7!}lX�U�ӟ�9+m5n0��{�D(7%�k�	�-�MY�Y0B��~Q��{�Z�Ѹ���	<wJ<Ƈ�Ԏ��`��櫺-E��Є��������O*�@�NR۲l��3d�5R�c�+�1�[����3��]��O+�S:�@�w1>	)p}�1%|4�?b_���N�4{�yV�+{���uכo����l��2`��aƅ$�����W�xWQ�i�l��+�G�uݻ�TƬ�;>�8���6���xEc1�i7�t-Q�����}W1��c�u(Br�ldNECښ,.$�"9-j=�
�������I{�i�zz�j���k|���_q��\(��}��SK�4چR�/�	 5�A|-� ���ᵫ�t��3=h���4��.u�<6դ���?���6����Csw�R\���?[��wr*zjm�P�\��_�✢��"��T�y7Dn��5kD$J:����/��1^P��@t��&�/tbFx��頥�|��b����^+
�����sG5Ȧ��28���cX@A0ȥ"�]O�+7	z��5�E��v$���x&��=�g� �W%���-y�Cx��+�,�+��Ù�G�bkm���V?n֨�)�	:�yIm�M����{#xz�.Z����6pc�����e;ֶE�	���p���P�j����<#a��gsh�o���>#�7$��)�ܳ�4ZU��Y*O�O8�7&�-e�TUa���]^^^XG
�y���f�s�R��<z|�21|��F���a�x��3|��'&�����@h����||e��xTχӴ��܆!���<��cC���H��4f�9H�}���so����s������&^�ѯ�`�7 �<9��v�Xf�R��ݥ�ۦ�&]�`y#Ͱ�
���4sM@v��M",>Q\���䡯���;�'a��]�+Q�&=x�/5��=[���P�t`wr�S���'���=�a���v�?�H��"(��]Y��(