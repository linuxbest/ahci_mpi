XlxV64EB    fa00    2db09��0�R�R��9<�� dzp_B�e،x�u�eu��oqԧ��&5py��8�al�[�>�]�8�b����r����S!TU'
oO�=M<����[�!)M��Ъ�AS�WQ<��,�e"k��֙\�45���hp��=����E %�Q��E��͌����F�Kq$C�Odqo$�2���ڕ��V��HEe���[-b?sD�Pr�H@y�w�B������3X �t���k���8����������WI�����G)�{�x����ƐL��X�z9ڟ��47���kE,��s��C\[B�":c3
�;� ��$u�|�鹔u��̭r6�_���5H�h|�⭬�w
�����%_�M�}�����YL���͵,Guy7cA����N�����J���,��)�q���j�7�BS ���������(B�P�+�>`e�e�v���x��O(��5�A�,-ь�%�u/�G�w�,�߶ÈX�����	� ��ʫ������FI.���V>X�`��9ao[����5ܟ���� �ꤳ���WP�y��9�T�G���Fuׅ�M�J��T���z#���� ޖ5�̦/�nY�S�<�Q'��ӝ�B�c���ޭln�)]�8+�LS�JԎ�X���T�F�<�J�@�͠�8,�i����؊�_赤�j��jE�6� ��=��x2��mI�%W��7�n��b�D��c��XI͛�'ޱ2��?�p�v������&�'��ノ����|`|C0&�f
eź��K���0]�䛘�~�A��%��Àx��J��3��a�|
}��@��	6G��JUi�m%^��1z����k1�܂����zz��r�gS_�y�n���C��\�]��l*���#��z�k�b|s4���t�%����%��#���O��H���z���rY��+�A�9NJtgī�,7(ֹ�t�(t$'H�liv�%"��RU��"�Z�`B����ѩ����h��g��N��� �r��0Vd#	���o�CSz�]���)����r4��ޏ���Q^U��p��FÀ"��K���%YH�kh��רF�x�X&��g�,ޫh�����G5��>
+O�;mr_wn��l���s�0��w�[�?$�=v@��/�L�4.qm��Q�9/m�>�r`xS��(Tj����TJ�qC�����������.��II����:�9�,�V���i����N�F�ke$~�4�W���e��R�kT̆u���*ٳ댕����U��L䟩T�.�||�v�9pe޼_i���)m��J�e9�8LE�͛�	#�:#�r�c�4��Ǫ�8�)����7<���B���$��졂a�~������$����B��N�,��˽�C|d�0K�m��^d
�hp�<���r:-������j�l��_�9j˒S�}���e�x�Rx{�=�l^�qN`�����37�K�T���(Zu؎O�3"0�iW�!]�;|kzs{�B�]B��x�)'���׶�%�M���dj��M�bNw����jT��]�c�� �*h;x?�e�����S&�v���O�R��2���[`�tC��.a�䴦�ۻ�����@�f�8�<*���?��ae����\o<��<����M6����� �B��V��>��(_���%s0=��Eg�U.s���FM�C�#�Ԧ=޿�������	���{�; D쯂O�#���4��Ef+
;����r��8b���*>�E��&�����C�>��-'��}�����i)<M�$P�U��C%�,����_N����%���Z9(����͟!�,e�fKQե�*�.i�fs��d��/4�����}��0��Un��
�S�|���9��Oh�U��0��j~�2���~!���8�����a3O��d;�0��]�(���yE�U��`؃���*J���v	j�2P�������z�ïT���y�=�EeL�������D-�h�:i�����G�(>o��p�
;��5ܺ�pEPB���:VGW���	���9�e.+�$��,�2c�Kk	��0A�|��CW��$�m�T�a�q�Z+��p�Մ��z�y;.���\�<M�֥1��t����(Y�ii�U�e���d,d8�{<L��*?�L�ר R'�Ds��H�T�c�<������e�<!ss�`X����%����`!�CW��P��I�ۿ�7�M���7���H�&$-�h��U�7�����n���>�w8�Ob^蹩�q�O+�vy	*� �!������J]�i���<9Jo�jЄ<����i���d�@@�*��M�#N�oO�ϡ����
o�4�)׺���4�@B㟴g~B�UX)��?�;U����I��\+�L%�����>"0�[��p���h"oU�Z4�
�t�q�m]�4�%��)��a�A���GR������)��i�߮�N���E$e�!Z���XV$� �/��h4$J����3g_�<#�U�J�S
���ǜ�6*q5 ���8�M��8��Gov�@<�ĎuJ�e��B9�F"��s���Z��{�b��ŏ�9Hw�vB���kO�+��,��(����6���Nf����\�[iI�ѳMں���w8���>?�Tq=�J��G)���l̞7��RT���;6�B���ܫ�X��}��D��ik��ƉV�A
e?�e}/�D1m�n�;g}Lw`�n�2��1�D�F�o�&�
k���#�Ĳ,����m���k����K����C�p�ǚ�ڴ^�ö��k��&H>��}�T����)f�P�t��ؘ���G���v�g�T�t�nuL~^*t�A�ӢD� !���,���cJ���?U̐f��g�	��+���N��v�ܨM�'�̹+��I�)=���5��;2G�M���G�g��1[����G��H�դ�X6w���*�N�Ҭ֬2���ׇ�\�Q���. �bx1� �S^�C���A�����dy�:v3�\!��k��|d(���º��W2M��M�8)��~vIGy�*{�k�����I�C�e[���r���JG=�y�_��>4߬��&։Q�7�]�JL�̽�p"�z�;x���f�ιf�(�
��r�>�����\J+t�&�������$\�*�����'�t���㾡��㽳&��f%�~����
SZY��B8dE4�T)���8Xj�>��
��|DI�/6��
�@�lz�X�;�/�9�Y�)��M�+睞@RɓI��+uU|�ÑK'�-� ��G<}G�M�:v�k�bL�k^��-�8Q#�Z7~�V���C�=ʡ�M[NM��:@[[�S2(��p�vB�o���Z��EЭ��v�r�x�c�WDeq��z�����Gu�-?G�~�4��X[_�mJӮ�$���f�OrTI��qcoo�ZV����4l���v��h�8��F����B�����ts� 7B�5b�V1<�����T�����E�X&(��n��#�������jc���ɡ^7���h;	:q�2hS JI�'��U�G���<ų����D��5LI:��IŪA��� �B��9�΂	UN���e��Uř{�0��Z�[�ac���3���Si���°7�������_c1@^��$P0(t���?D���9�İ�����z�B4�!��4~�t����r\��vcI���~pX��a�y(�ȿWH[�]H�=��=������{�#$���4�h��x�i� }̈́�>�Έ�2Ұ,MJ�"O'5C��L�4���D��m��K��*�!>�+���3�5�O������KU���iy��wu�cxǑ�e����#�eD �9�n���I�:�Ky��&T�򥏡�h��V��y�L�{RD��@:Ϻ����e-�??�4 0��N!B��s�f"9g���cf�*�9�l��cwxW�����Q��y>�+
{�z�OAMsr%c�$��Ԫn�� �ߜ6l��\��`�=&S���|(o� ����b��Ґ��(xC�<�D�Au\�*[���V��R�#!���ݥ3�D��:]�lm�p*�O��cJ�������/�l?<C������i"�7��������m�h��p��JХ�G��C�C��c�Y�mu�0�L���/�@��6��3�䏋)�D�����=|>�#�@o[O�xI�/�y�5+�y�qre3:�:E���B�{��1���N]�I�谻Խ�>������Z�U��#�c�%1�ޏ�VU��Cv��1��)���1��0�Wv�9��4�#�MwMu҃1{O#V�~an�A�WR3���e�>3C��|������tu��d�茜�����nh�B���R��,2����ē�P��5�W6Ÿ�H/ҿ��9�0�gC�>f���^���g��O��Y�Y侫\h�`9 ���҄S̠ɥmv��Î���I�8��r ��>(M_�|�tg���DR�e�����S_���G9*�Ϋ��?s7����/�i\]ݕ_�
{V�/��K[����?޹��}vF��]ɔ6����(l�:l�$/�@]y= �/P#�Y,4Α[��nS����t���	%���Y�S���[��&�!f�X�W+�\�-iȘ\ ������w��@9Py���0K�ӂO	�NH��)�ꄰ�)���Ŕ Idr�a�g��EeF�k�U~O�"�M����A�C�%�ś(�4T	p^�]�Ӿ,�Y�@��EU'i'�F���TM�qYDo��^�Hu@�b��L�;ݎfX�ܩ��,+��>
_�h\���r���"��4����Nv���_V�aE?(�U��!-I�}��Vl���V$�������;<fO3EJI��Po��J��[g�^&��?���J�U;t������̬�����\��k�9�)J~K& ���� RzS1����'�0�/��F�q^��� 1^�ʹ8
I�ꔢO�ø<�t,����f2�$~sca�B��%?c��s�*}mGi����I�o��ڰf�M �
^�0@vw�~8I�9�C| �5�iv1�Ux���>��f��b&�b��극Վ����okȖ�K�����������U �y����P%I�Gl���T]�p�+�Rtx�:6�)�k��0,������G){�%7���z��-Omyȁ��q	ώ��k������'�eq��t �ь^q�~�j_�\�V���R��i� D�ZZ7�SP;��� �ǭ�n�;�g=�z_D>�cN8�h#���?�����(��Q���V�0�Q�ɋ�{@������h!>N�w�����|��N�ܬ���+�mW+��R��)#���V%�>��i�O���̳tk��Q�͖X�7��*`�7ץ��eg����r��Ʃ<�kw[wYOe0'O��)kη���3��Ա?�r�˩=�B�Ug�(��=�ʇ��9.+��|�۹
 �ɷ7����J��f����i �^���a�:�tl:\�S�D��b�j�������<
�P��z��G�Bqq�=U��P�Π��4F��b�H�c��or��I� +<�q���7��O��AS�n'��� U��.�F�Q�������B�fT}�6�g#F*)!n�B�c�A�.��%B���W��f!�<��������D��u�"�K��n��j!�X+��4�y~Aį�"-��^2%���+�1R��[�C���;3?�����L�c�$�1��"�DWq�
&���n�˔��Qg#��^�o�۹�&d � �ڽ2/����+ܠ�3Yi���f �F�[��#Y;���mԤ�7��S���/��ƃ�UZ���#�'�%�,����X������2K
�c�E����ͪ;(�,F�oa�(��I��?�2�$mr��B[�+���f5���T��ly��ȭ�rZZP^猘t|��,�#�Uxr�B�aѺN��UEx>/� �9,�?�/}ϭ�l&5��N�	�B ��>q!`?ݏ��&"�O���±
�������~��/����3��S�AF'{�{T@�?L�bU�,�D|�/IVu�ƾ�cj�6hӤ!I����+�J���xJw#k���iCk�X@�m���g��D,`@g���ڸW���:���&����������N;���E֥~�w���f0ƥ���������u�ґ�g'�6���z�i�Y��b�Q���{����k��a+��֠= L����r}�'-� �۸ �tz�dؽ9�f�(HJ"j5X��?���� �����^�4����x��U	V�QA�N�ϩ�w��I�i��В"5��-�"db��I�����=�L뇟)���!��MH�#փ����8�mr��¬��;hL#��ϵ�fv�5~!�6W�#>�F��p6�A:K� z(���1n5;[ȟ���iȬ���6�W���
��Uim��`ߙ�֋�%�jNߕ������jq����T/��
���q�7��.�����h��ƞU	v�o���M ����Ba��ˁ1�}q���nriVZ��r���X{�!����n�h�*�-�(t��%5J]Md�i8�?mCJ����FЉ������[9�ko?�����bh�G<y�`�5���KyH+)�O5#�c_��Uf
��"�F5�\�s或�$ۓCt6����#�;E\���:��?��گ��vQ' �;����D-���H��EW�Ϯy�G�Ł��3�n#딆�~�;���'�q 7��������v�Ja�X�dtމl����JtB�#�Mm�)�L��>��AQ�vW��ˍ��me��\����,̐@*�0�,�d�����K������|e4����'p��[|\m�Xn��k�fd�,-g���Z�_m�7�S�7ͬ��k��0��m\��p�3�����$�˷�*?�#�y���>�%��=л�촧1ܛ�3kg�a��:j�O��nI�Q��^A�s���3�kV��8n��j��LMd2��}��-�x9���� �\�|,����w�����$yD�� B��w��̯�4wC�V�&��hϠ=�@��gB��+4�8�:Z��*��e��}�½ke����B!���_:>	~Q	��u��4����x������j����=S@	�Z����7�ٞI���7�/�f%���x�cn�^DAP`5C�<�\=q��h�agZFw�[��`y�M��tB�8�ԑ�j����"I�C����RNK�(�8��u)>$�k��U�]	����=�rNw�e�h+�g������"+�5�.}D�K �:4�5�Ā�G5�rgV��wŭC\O��DWm�u�<��{��қ����4����V+�x�q��2y��oW�kBܝ�+�K�=`���QR���o��ߩ-��j��:/ԟ��4}�b��?�PC�GGާx��{`C��~�+EW����L� uE��
���#u�Q���l��o���� �F}"�J�@����=KJ�L~͐����_����O�6^���ZR��u9��H��@�I�'�Yoy���q��2��bZ�J��.Tc�rh㰗�\��@���Xp�[Q��CZ����ZxPɩv*�=���s9�A0.��ȉ'�-��6Aom�r:�k�3̇�#X�#G�Xdo&N�� ��)[
�)�Y�M�����t�VX?�٫Eț�)ݜ�=#�>ί{��_�����j?�O��/��R�ܖ�	m�4t/������l�평���&7��E&������X��n8������y�G�B�j�����\���;�6�m�T��E��3@Ϫ�K���8�W��ϔ���C�?w���E*[r)�.�����*�aL$��oi�G~�/��@;�
��u��T������C�$-oR3ɐ:��%��4�y`��w���L�&On��_7��{��Y!C�n-|�B���)�'����R%�ۜ�؜��d��^�r�`��#�qfUX00�L��ΤD�B�w�w��+� i��g'����!�3�-?�VD��k�O�Wh��Y֡.`���D!ǅ| 𗨽r=�*/r��9B���de�ﭧ��P�?	��W+��n��j>S�d87i��^���U�ѷv}w^q��W��5�?�IKrb�?X넲��Ck��Ʌ1>R�mD��'�W�y�bz��a[��]�xW]C:/���*5)��ZHc���ܝ$5�Q\u�z�0��//�m�Ҕ�ۅ�nwz�S��.$�k���֦b��MI^r����B�C~A�N����E�:ˤ˼�?ԏr�F}`9/�+��$P58E幱7P�n|����{��@ ����h�#S�K@S��r�s Is�V����Sʅ�T�D����������@u{M:I���U���9��׎�Kȷ��p����#-�W�u�4��������|j�����r^�C�I|��Mg]T�ŴbqOzQ|��#�Qc:�>*�<C�D_�&����ww{�9��?���n�M�8�������DĲ�d�Hz��@)�j��~�nucr�F#�8�0H^p�P,2V�f��qB�ç�L���ks�����kT���������?�05J���P������y�UA+��ZLanC5�ȃM�F)���7�!���BϽ�J��=�V��U��./���2f������,��a���N�M�ޒ��·-�d�3D`~=���S��m4��L�Ot_����Ѥ/�<n��Y����rI���B{@e|�S
�Af`�.]X�yE4]��񃌖�U�i�aR7���<�s�����l�oR����=2_����?�zXM�� V/�� t�l
f[�xgv2�
],�S�@W��'G@M�!�B����oA��*���1Ƹ�]����+��1S�p�spD'� ���@���2�լ���]0�h^�IA6�oN���3|����Ç���IM5���&���	��D��%g��㱈2'�<;2�OF��xCæ�k�@9���R�Ķ�˥�p��t
��AjD�X<��e�Q��-m�( o c�\j<�.8�a��;�
1��j�b���s����*���{y|����w����n"��Ε��:�)\ȧ��XI�K6-�Nm�:�?�'�{�Â,�`��T�\a=�۳�Z���������c�KR-��yV����ۆ�� �%p-�ڃ�7nvm�5����Q(��|L���;�h�q4j��t�9��8@�|k�=�[7n1 ��N���e$�H�3Ş�V97|�\ qV���ڧh'k�\X����KWJ��ՇO�ځ��s�	�$t��[��)q#���G�1?&� �~����������g]��̝I��@Q�O,t�fƹ^&�h�x&&A���!8H��i���[)������"�����>�bk)��N#G��q{֚J�9	�ؽ��Ϫ� �9Q�!�(����P���ZuVG8���I�4��y��,t!@ ^3���P�����@H�=3�D�ru���`���r��M(���~��)z)|m�E%��S���I�j�R�[�n����}��`x[�l�wU᨜��Ř�$���*�Ѷ �A�ɬS��ӯ��K�hu��&�,����[�z�0�����.��f(}1A��`OZ
%�Z2A^g��E��)Q�*�U6�k�
�O��}�6��ۋ��������b�o��T�C{2ȓ� �O�hщ��
�#m?^��+ԏ^>���'NmHYUaV�E�#�3�kݴ�H����x�(�U2rM�ç�T`��,���vP<uT�zK�=���x�4d�U����<��}�{�/׃V�Z�jԀ�g�p��������g��BHBⲵt%KQt&w���1y��rX)�V)��+���_���a�m���Fq�eve 5��b�2�u�5ض��#�,�C��|[���>�|].��;�!{Q���~��8Ҥ���1�g�l#)&���8[!/`Q@b��lD�2�ƺ_��~q�Qe�
��g+a���QP�";e����)=�:VS����b�#0n��7���Z9Ԁ�څ!<_�sbd4*~U�V�#��^a��5�1�!y#Z�x짠��QH���y�q���]���2F�~l�����b]���4�����p��d��՝Z�4��x\��@��G���fͬ�|V��F8�Ȉa��o"�~~��Ѵ��-���Q�>�(��w���],���v�B�"��%js�t`$�S��╏&޵k�O.�����Ŝ\Aԋ�_=��OJp�BDF���9�/R�R����(�����)ҸO����?���xyh:d��?���K2�LYQ�k��o@�3�>��D���ت�"#A��?��4�d�	:�v��Ϙ��V��|Z�ʼ�8��5o�� ��˷�߉+��"���*v�\t��P>����,TE)SI���t�让���:�9qK"�ȯ��d&0K����������)`k��`�ʦ�y�H��qAC�zY�ݰ;<��v>[��%3fEK@�)*�����GȐ�ڋ��F�U�-�P�	Ak~�`�\Pt�`
�f��Cs�
�%E�����)��QWO�x�r���4Z?丯ђ�!�֚��A%�#{a�}��m��F����)�+�ˈ�jj�7��-�ϖ�7����[�k:(�P�9Cqݧz�l����Bz�a����V��a��TnH� 4.�]��N2���z�a#���P�̞�7�E��p2�jw�n�Q���#�^!x^ B��@��� M�]����03�@��b7�H<�:�&�*�`Cҵ���X>�m�+ǅ��h^ȱr[g"����	$�-ؓmR��s2�s��T�a�%:P�j�@9�1��}49���M���	R��2���#!O}6Kɼ�N�}�L�� �[ٰ_��WLe@]��8���kU���0����"y������&���L�L�_i1;7����1��Ȃ�XҼu2��-���Ud�22��>�F�)� �j���_�V2�i��Z=�tFN�ߖe��t���
�ɾb�uX��H�j��hۏg�`}�{�<�}�Ľ��|�M�b��̩F�.���.x����Jl���}���b�[��N���J�͹?uإ���ܓ��g6�w�I�@_�$���'�_���^��C2�Z���&ex���6�G����e���)|����V�{�)6����e9Ԧ��!|����7a7�h5�n�[vb��P��f���*������smV��-����{�D��S�� �7���q&�4���Ӳ����X�Z�h!��nmў�/>^&��4M<� T\C��ȍ�Q@(|���ɒ ��l|�!=��'xV1O*� �WG���iD���dߒ��?c-�6@��-Y}0++0�,�vN��:�8U��S_U�B�^��3�ȩz�J�h�u�;o�wXlxV64EB    593a     df0>VcY]��W��s2�S�C�^����"�rF�jݐ��քvd���=�D�{U#���3?q�V��d�pK7 ��|�~�'Ŭ�s\�R��Ё��\7����$��+n��L��O�.����[�=��RXjv�)�^�5���r;�0�i��t`�63�z�v�=�;)���"�}oG���ڛ�u��@�ANiZ.�����	�oZ髱y�Z� ��~,�I�+�����g�Õ�L�C"	���*#dJl!j��Z �2 +m����_������;#�C�k�R��Kg�].��t���f�ޱ�%�^N�e���'｜�D}6�jޗ��߳#�U���(��3d@Ȥ�]��;�y%��MΝ�� j��`Ė����ș<�l����!g�����ac/���Չ1[��z6�������Ǘ̴�/�i��3G ���~�h��n�e�J���81��Pf�U�M��1���oں䍁���VzpJ�ΪҦ0D����v����M.���\�凍�;ۘ�=Eʈ����iW�%�g��<�Iy,d�Y�[�k�e�ೄJ��y��uOQvz�q�i�^F�@K�����#enf�y'��"��P���$�͐cg�����8s��غ����i_���n���]%*8�;���
l���6G�|�M��Ͼ�l(��`F�����4�l�u�YT˳�vg��Q���
�p(�#~�d����&��Q�?�
��M�[l3�W/��6=�~�E1YD~֔IZ�j�q�q�e��z�9Q�6,G낅 ��R[ԣ\�|/TҘ�ϔq�:�?�P�%T�Z"�����y�N����5����$d{�*JqƺFm�@��(U5�	P�k'T'%YX)!h}�3к�����o�л��0�Y�Tg\���W������mzݖޘ��#z���[pҺm���\
����ܔ�;?�˴�y�뫠���x�L��I�G��?K��#,��!c6���U��'Q�A{�� �֝�8����B��]8����S�2���7Q�/�c���v�.3�Fk��$��S�܀�|�3P���en�5�x∑�nOX�_��5���*��%�^�����f��`�+��T�� ��d��h�v�2~MGL���V���ÃSa@YG6��U�@�Š^0�U�c�˸u����	;����fP���X��N�R���:��oB~��`��l՟��<+�I����h�w,M�1��+����G���W3`�����|�xQk��|&c�ь���q�H�{K�DF�<�R�/E=4m� �e=���n	Ǳ�.�S!/���v�|�!�G�U�Z;xD9H�2n�ߘm��#3X��;9~cY�e^SC�ܑLj����)��(i> d��B�9��
��LV�
}�(�b���z�i�,�k=�Ě�	��!Y�;~R�՜�kE���;��U��0$��?OG�c��7�,ӳ���Y~�ɔ%5�:�Uo�=��p��5�ɯB؉��	VY)�ͯ\�j�c�wZ��V����IPȴbX:8��_HI:bFy���y�4]��]�ό$�v�''�s�M}Ƨ�Bm�v�
�|�ou����
0u�aV�w#+��.�<6�tfT@��$X�? k �x3��)`�,y?e_�O�,$�X�hg�)-�^����z�8zky
��
� L�?~�W;��lbWx8h�տn�<�E���������1���[��ӔW&
�ܸ9���?6P�ZZ3R+M��bod�����ƱQ 'D��C�M�`yx�9�>Ͽ�H���/�S�� ���(Q6ذ2=�Q� �V��l�U��7x8V�ZZ���
I³���&6��f.b08��w���7)��4�Z�S�Ei��L�x5ԃ�b��%��ũ.7��k	 C��&
޶��k�Bfh�[���>���o+�wH�xҒ�"�������P{lPةhe��;�J��#X�tIV����Xv'��1X]��5�ͨ�DVI�.?c/.4���d�t�?6�ͨ��K ��z�F�Q\!]!2��gg����Tax��F��?�1�,��������.�l��}�fz��PL�_�G��+X�<|tf�r$�:�҄a�����T�7�E�H6���d��["�W����P�b�<A��@������+
6�̽�b��s��9�{��z���RU�N�Q�����?^{[{�W|�5��mdh��[W���f���d�F����<�z4�[[>����uI`E��? ��k����p�F��K��E��%-���kNƚ�]U�ۥ`��%+H/L�����SRQլ7L�1}O�70	�LR��-�\��}�]g�Κ�yX�s�a�9�Z�ZLxKa�̏�I�*���H�p������$�2��' �en3a�
ֱ�er'�?���B\�
�R�'O��uԞX�֟3>���Fo�F��|*�$o�������3;[��Θ6�Q��������a`��m<?v@'���,�jW(��\�soa�Z��}��3��M�苄�;�Ԏ��-�c�l�Ҳ����-J��{J������uX��6�����M�?*P^J���}��:�%s�}�Y���@h|�×�$����P�?u�I<�4��NE	 7���v j��Aj����t{��,��Xx̽��Q��v8<ިRQŰs�8,�����ș-��k�ɈTr���	̡bC�i��{��#�����h�K�fm;VѼ�ie�6D�������z�������;^4�^8@� V�L��r���oi�$�*3b!k��P+�9ü	��i��Ɏ媎'��H�(�9d�U�Xsh�u4�����U�u�:�R^IߒV.���=�XdSi��V���b�D�����U�g���/�Ɖ+�7�J9�>���?��y�2@Wd��&l�=<��O���hE�
��`����,�� V�K!�q���ϒf����#�R��W|�������W��=4/4z4�񚳰aB�����@�֞���,2��]`E�t�n����aLǷ��Τ�u��C~Zqe�贚�`��jDO]��P'���'�ĳR�;%P��4��7ڿ��6H��B�%/��x�x
���Ҵቍ"0��s�M4�F��M�/�8g�؟ϐ� Jĝ�;��i嘵���K�,��Y��H��Z��ږ,]�uj$�LM���x��Oݪ@��Mx����/pXJ���#j[�m[�
���P ��E�~R_ʳ�}���0V��Q?+8n˘�8��s����_Wa�9��O���z�Q8k�W$j�����B%�$�y�SV����ۯu�m�I�S`V��� �7�2�s	����m>��6hP���ϗ��b�HWR�1�D�U�/utP�{�flq@�=[=�i�Y�����+5���I�@?3��&����Vi;�!��#܉��QOW���d*p�f�)���#�����Ah��Vn����`�#��3!R�n�S�Rb��D�q8�҆o�D�l�4}V揍�`.�1m�#��K�p͎O��o�,�;�y��$?