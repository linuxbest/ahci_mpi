///////////////////////////////////////////////////////////////////////////////
//$Date: 2007/08/01 23:10:49 $
//$RCSfile: mgt_usrclk_source_dcm.ejava,v $
//$Revision: 1.1.2.1 $
///////////////////////////////////////////////////////////////////////////////
//   __  __ 
//  /   /\/   / 
// /__/  \   /    Vendor: Xilinx 
// \   \   \/     Version : 1.7
//  \   \         Application : GTP Wizard 
//  /   /         Filename : mgt_usrclk_source.v
// /__/   /\      Timestamp : 02/08/2005 09:12:43
// \   \  /  \ 
//  \__\/\__\ 
//
//
// Module MGT_USRCLK_SOURCE (for use with GTP Transceivers)
// Generated by Xilinx GTP Wizard

`timescale 1ns / 1ps

//***********************************Entity Declaration*******************************
module MGT_USRCLK_SOURCE #
(
    parameter FREQUENCY_MODE   = "LOW",
    parameter PERFORMANCE_MODE = "MAX_SPEED"
)
(
    DIV1_OUT,  
    DIV2_OUT,
    clkdv_i,
    DCM_LOCKED_OUT,
    CLK_IN,  
    DCM_RESET_IN

);

`define DLY #1


//*********************************** Port Declaration *******************************

    output          DIV1_OUT;
    output          DIV2_OUT;
    output          DCM_LOCKED_OUT;
    output          clkdv_i;
    input           CLK_IN;
    input           DCM_RESET_IN;

//*********************************Wire Declarations**********************************

    wire    [15:0]  not_connected_i;
    wire            clkfb_i;
  //  wire            clkdv_i;
    wire            clk0_i;
    wire            clk_2x;
    wire            dcm_clk2x;

//*********************************** Beginning of Code *******************************


    // Instantiate a DCM module to divide the reference clock.
    DCM_BASE #
    (
        .CLKDV_DIVIDE               (2.0),
        //.CLKIN_PERIOD          (6.666),
       // .DLL_FREQUENCY_MODE    ("HIGH"),
//        .DUTY_CYCLE_CORRECTION ("TRUE"),
//        .FACTORY_JF            (16'hF0F0)
//      .DFS_FREQUENCY_MODE         ("LOW"), 
       .DLL_FREQUENCY_MODE         (FREQUENCY_MODE),
	.DCM_PERFORMANCE_MODE       (PERFORMANCE_MODE)
    )
    clock_divider_i
    (
        .CLK0                       (clk0_i),
        .CLK180                     (not_connected_i[0]),
        .CLK270                     (not_connected_i[1]),
        .CLK2X                      (dcm_clk2x),
        .CLK2X180                   (not_connected_i[3]),
        .CLK90                      (not_connected_i[4]),
        .CLKDV                      (clkdv_i),
        .CLKFX                      (not_connected_i[5]),
        .CLKFX180                   (not_connected_i[6]),
        .LOCKED                     (DCM_LOCKED_OUT),
        .CLKFB                      (clkfb_i),
        .CLKIN                      (CLK_IN),
        .RST                        (DCM_RESET_IN)
    );

    
    BUFG dcm_1x_bufg_i
    (
        .I                          (clk0_i),
        .O                          (clkfb_i)
    );
    BUFG dcm_2x_bufg_i
    (
        .I                          (dcm_clk2x),
        .O                          (clk_2x)
    );

    assign  DIV1_OUT  =   clk_2x;
    assign  DIV2_OUT  =   clkfb_i;

//    BUFG dcm_div2_bufg_i
//    (
//        .I                          (clkdv_i),
//        .O                          (DIV2_OUT)
//    );


endmodule

