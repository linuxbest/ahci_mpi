XlxV64EB    7a1f    1a20R�)�<��55ɯ�aJ���ڟ0�#��r����XYK)<����u����>��\	�ϣ����3WÙ??3�^Y� #�l�:IA̔�KV�a0����9�e�9�[�#�-�1�d�`��|���l޹�Y-�a���X!7�(-by?��F���lv�\��Z������Z,�ΩKF��7�H��d���j!���P\%�ZVX�it�G{�F��\ W%�C(21�ϦH�f&*�o*1ǫ�Jm�N	���a��W��&�R�%�S��o�$f�J�Aږڈ��W�P���1�q��ղ=���,[%x�R�oԨ��,�
S���l�
��h��eC���S�P,V�> n���j�2*�-���̼����Q3]JL�
V/�?��b��۱g}�b9�>7���@��|љC4L���gc��v�.�����Ȩ�N�|�d1�x�{Z���i�v�����F>[�y�����z�\�������K1V�ɑM�ʠ�J#�Z�uz�ޕX.:�m�5�D�g5��!`Mf�#=ն�*BG��y��	JlR������i<I��Z��зz�G90]i@ͭ��d؋�d��x]݅��@58�6���S�h]������)ȳ�)*���"ٯ%ex�g�Yc�������%�9T$�/b�� _����Ʒ��T�J���N�r����H�4�e�(��j�XH14Xw���I�M�u�P�q�E�V���h�r׍�4!�h�԰��ߙ`�I��`��+��=�P�}��6�Q.5�CFQ��Sw��Ʀ9��ZI�wy�6�J~AF�Bty���/2qd�x�䧺��Z� u�� K��~���( ����
�'�%#[ LA�l*f!s뷥���-��G��rBb��5 �c�1:��z���|�8�M�����l@Ο���ӓSo\2���B��D��x0�Bs�ř����!�d+R��
�b��vxD��~/E�������}�bc�F�d�_YP|cÌW�r�)Ui�z?��\7�u���{�.[�+q�_.�\�y����32\c[K]��J?I��eD[�P�#J�E��g� R �$7$��y�nD���=�m<@��M���H_[�w�i�*�݊?�f�J.�]��\lY4���n�\פ�W0��=�@j��]�Ĳ�1�
�%���쳖V6���u���
��5a�]XE+
����Z�<'�&�7����lNGBc���Ӆ�T���țUj&#��K�O���_�x�0�{��~CS���7�阓  ��u_c@�:�,��҆�V �?�����|Uj��<��ha�E)�,%4���Au��,�R�k�lѪ�7������ K�˞���a�}gÀX���`?<G�m�:MKIW��:��H/��@x.��
��36�t���B�W[j�$���Y�za�M��=���)���'���<y.!Qh��x��%�X��l��'7��7�'��?����_��#8a8���R s��Z�{j�z��䪸 ?%����v�,��L�-�&�w�ϫ����}�$͟�0�S�ʁ��!7�z� a�@�<	6$;ߒ1�� ��Kw�'�B�Z^�0񓢓������/ە�0�r�����7��mFz�Ͱ��H����(�w����֔��wA��0�0�ֹ��8��1-��'���	H��f�!��l�W��
�B^��V��fq�Q)>��\�t��D�ǔ�ߑ×��X��ἡKξ�|����`	�u�5 �#�$Fa�O�)�x_/}!�����o�Oj�9@_��u��}\F�vu��ލg�n���
����mSW��nbky��E�:_p��_�
6Ri�����{�h�dvx1�lpل�!*p���s���T�'	}J�aQ�̼;D5d!$��r�n��<:i���֥%�gi�2��s�6�Lݝ2����@���ĕʒ��p� �g���AG��;lቬ|�B�����b�p��F�De�ajY�Y�bc�w��>�m^���Iɣk_Qg����O;��>e> �>뼯��'�{��5r�����HL��G^3��C�ś5�7(�L��w�p�=��h����@D~W��] �6�8��7���1�|�3�^[�� w
��3N�o,��g��s�d�6ΖA��;� A��8=~.Pt.%t+��Y)��xԑt.�Q�S��\�Rn�� pW?��|�Ø��IM��p�Io����:�g�� ���T����/�\����0e͇�Q�=Ŝ�_�A�*/3H�,�q�|WzcD��pZz,PS�A��|��)W����冐%�܂�d��Z�\f��W�Bg%���k��p�`��PS8z���z��Ub�(��"��X:���	L:�e��X���(���!�`h�򫇋#�=��k�1�Z	�[�@�u ��GN|�b�Z��V1	,�J̜��z�F���M����a&�4n6̷��0<�m.��>���̑_�D�k�����&ԃ}�辅bF&%�x'-�
}}�Zd�r�{Ys6`u�-��Lk�	�� ��D���p9���V�e���!��kZW�=��-�= ˴�L�*~�!n�v��~�.���m�Pt*��f��(/H<��;]�:�
|��X�P���]��ae����낼0��eW,���KQ�t�~�ə��E��׌B��6+�U��+��Mr��a�_���%k�}H��S{O
��6OSOG���1`������l����"#�BE�������XC�(Q!UM.�f�hS
]�uю5�_gir���[�$?��b�9��vB���?��]�Z"����)gT8	h�jx;���Lڍ�r�*�9s^��a湴$�'�G\�2�;�h��BJt�.㗔���r�D|<�������p��e׳�� m���̣��y	�QY�6�
�	����w��ÇU_�C��76��B �|�<c���g�Ge���&�� �!�Zb�I�`泧~�ة�&�
��>�ڳ��b|RД �b��u���|⵺��ͿE|+�}/Z1��{ �К��nݚ����aʂޡDr"��A�,��C���;���g�� 3ϳ�퍔C��ub�Λж����G��<�H���q �D��|���h�DqC�9i$Lp*W1ŕ0$�[�$��H�.s�"�U�RD��Tpu�����z��d���ݥ��*����{�t �	"I�aa�wn�cz�*M��f��Y�N/�-�UV+��J�J�Z�*�������xn1M��]����!'�3c��`V�7�(�4�V0��>��s�+.)�,Y�R��!OTI:A���+�%lp���`��=���������.���R6A�4K���GvҾ|���tnYer�!�ʇO�����y�:!@�� �E�2�=Cx��"�A�踽���Q��
��6$�3t�Cq��)6����j�"k�ז�w��&����t`�4�:�|%�u�����7(��qUC�&�k��W܀�m5������KF<������cpG4�����Rk!�,}��1�9�ҥ��jN���Of�{ N��u$N�����'�0d%#u�*#�=Ȁ�d[,Yd��T���&��o�g/�@�$�>����@7o�=d+pk��)����5rV5z��݆4Y�*��H+Ez��"ф���r�}�z���k)Ӵ�O�PV�c�����Y�&���&lF�P�k�3W�d� H�
�]A�˛�b|�1�3�u��)��S�x-�r}�S*3���D.��t�����N�Io�]i��F�c18���++���#�a_���%�꾜��(�V�zAN�+�2h(qs��c�_�����R�][|��\;�	/-e�]Mo�t�u���1[3�CX�"ҔP�9����ˀjt���<����A��26J|{�J0�81Zԕ#�����`~�kI���'߂㳿�Z��:����4���&f_ˋ����VC#));��*�{	Em��w��t5Jӝ1�Ch�t�"�]&l� /�5P���u�<3�����R�?�V�(��,I�C��O�A\Z
Z/�i���/q���;����d)��)j���9�dʋ/ڜCQ�)v2��:�G�O�l^J��[�$����`�F��Ur�?�'����K9���m-���7��a��aU=_��Q���7(�1���Ha�ATn����d�C>� �#t�����x��^����S���;�|0#F�G;b�_)�hDtA��R�As&�:��YP�v��s<U3��9�]�QY�%�������T�Ao�-�� ���z��Sb��6�NM|��P�S�V��*Cx�O�!-'��󧗬������� �G+�▅��zȗd?T�A�.�D���)�M�z�3��׍�*ʪW��[�0����~<[�T�:== �_�����(O�o��z��	���p|�y�j&���HF6��k��X�!�l�kH�N��9�ݫt��.-��{n�k�q(:� �t�!v!翭�8��S���N�0���f��n���(,�F��/o�M��f�S��餤�GK� ���8�n�^3t�f+�m@M�X�b�]-��&�Ν|n����XEW��=�.1Y8��Y�Cz9����2K=���Dq@�7x���s�LU����kE5
���s/��N��ct��H�3��E+�5bz7ĩ��Z�>%��o:.-zZ�n/��X�S/R`+NTN�Y(Ze����B�:~^*����i�@���ŽԔv�B���%GΛO�Tg�*���*���,X�v�{�R�U
�r�I���|hk������Z�	�������	4?�(�:^�T��*st/\�?1�ݎ~�2�e�xno��ȗV'�����4ZK�C����G`��\��3̪�}(�)�jfl.������az1��=�b�6�ӻ�Dt�k�l��<�\���ǈF�R���yl�;v��Fqؙ� 8"��x��<U���E���X?�d$;�j�����y���E�:M{~9���dY[S�K��8�GE��k�N,y9(����<�O@p���M괹��kn�bʍǆ䞁$~8:�6{��Lr�;�3{�ݓE".�tFb��-�3�'�����6�,<�_���r�"$e˴f�� �a�U��1!�������(<���Eܱ�~�[� ƃ��u��]����IGTT2�'��u
��V�'ޭ<��Uɣ�h�|��D������'�9�3��`�j�o����	�#w
�+�ص�����o��bw�T���
_��1D�LQ��]�'h��~t�/�G��j�
��5�5ڔ��c���6�
H�F��߭h0M����M[��Z�k��J��݆��
l�3���;5$���Tm}��ٯ��iT�^������i���h%�L�=oG�.���U^�K��ȧ��A�!'�d�^9`0�%�:ʹ�b���+�/��QG }�6�J�O�d�6F� Ǹ�3��K��w�-138��6�l���5���m8��.��C0`�M�]���4�UMH#c�0�EǢ��Kf�
���#�B� ?�:".YjU�e4�x�k��*�"�-��ݮ� !�}� �U.C�ou��;��⿡����.±�P�,���d��J6TJm3f��~m�����X�d�1l_Z=ϯc�����Mi� �Kx\�r* A�H�ψ#���!:j.�&B�R���}�R���AJ0��b����c ������&��܏� �O��S�B4`��D^��[�~A�m����!�iR�s�<Nt����Mh&�dY���ׁ��:�@cWN>�\t�4��|jܼ�CS4mH8J�;k�c͘I��Sy?qW\O�.rJa��$��]�x4��3����D>���m�W�!�k���=�L�e�2�}�'Eɋ֚�@�eo.�
��l���6��R��74�1�gT�ˑ@u�,��kMX[EA]e�Mk�w{)O6`���1��÷���}�}7ɀ|g1h �����R�N_�'e��+��";�4?��[|��/�!�
�^�h�)�������sd�YV���%�Y������0�\`�T�4�I�tѨ_�84�3p)<-cP˚*Tlq�V_d\˓8�n�+[9L^��F�joj!L�f�^'�miD"՜O��@Y��������ɱ[;��8�*"[��UY֑\�A���i�l��CD���FI���?
�$p�)�������<L?��
	P�=��dM8����d�L�>B<m����:�p�0
S�Z%�'mb���Y�A��i���S�,,\�B��F�	ƥG�ܵ:䤵����#��\����Q��CnV��!#�l+���d�,.@^��Q44����W��iUG�7OW-�u�[:=(�����n��LWz��Xi(?��f�:�:[����p1��� �y��d�H nP�x	�)υ��@[׃JƦ�p���Y�`k���7��z��i䑤�t鴾b��W>���Rd�`�"�,�	���x�
S�r��gn.q] R9�����:S@YT���Gl�d�AJ��K�(�7�����4�͉{i����yR�)P>���F�Iu`׊����P�C<�1X(�V�� �M�R<��������