XlxV64EB    59ce    1410W`���Z��J�g��J��ԣ�
hC��zZ����e��p��0�� N�CW���PȯD &̉#���3������9�CE����X�Lݐ�%�3�1~m�	���?!��frg=�sr����uip�y�������S=g�(R~a��8I��$�#��K���ø���X�T!�P]�U�5pg߫&�o]�=0��.&�A\����w��_�ˊ�)�Ct��²�I��7����AD�d'R�&����R� �vb����xں�
�u�C)�5U� "���^aS��CD���e�z�b�7I'�G�4��l<�W?�[�����kt	۟�:�wJި˛��������bV��rH	�o��A�C�WX�����Q��j4����I���IdŬ�jz9�ۛ�K�&ܺ��l�� ���u��������Q���xP�S�RH-���HP�3�f��ϰ�F�����(�iz��1�5%:@	�>
-����<M	&���?� �?C`��=�@���ŊU�Ŵݞ���na���߼o��TYZ��a�+��
' �G��X��h"�"k���W�K���+�yt��O{$Mn�}e�vӿ�PI#Iܽ?�Y�W�����N"���z��9'�U�WD-t�l�ν�q��40��v?W�K0��)�B����E�	ªR�n��Wo���p����L���q[WEqNZ<":�	D �e�F�j>�}����ALp\�AC1���٭;�\�CRU�v2>�t]��m�2Xf����|H7M�.��o~��z;n#���E��bB0RMI��&���w YD�7+-& �_X
J�z������(��"Lܑ�䭒" A��3�l;[��(!A��\6F��`��鰓�}1OE�vQ刷�F";v��1x霘��� zkxDJ;/����e����؀dM�����?7y�s���%��]�.�c��\�g���8չ��`� �sQe���V���h_��b�X����k��4���|x6m�����8�]�sM���eZ����� #����.|割r����+��-/M4����TB����sE�^���~y�G���*&��u�wCǱ6c�}UP2��ӾŪ��jS�M凃��G7�֘UP�J>����ȏ4>�C=�M�j����+��Hu��'
���#D�1(pr��O-ELh���;s18t��A � �,��ܒYn+ps����.�;1�f�G�+�1{�x��<r��v>�8��
Hea!l`A�Eؒ�-#5��no:�v�^;��9� %y�h�O�����޻Eb���p%p(�x]�?�k�Æ��{>��8���f���s�N��_/�L�tY'ǝ�"/�*@n��a u;&���+Y���a��Fb�4�������+�>������7�`ux߼�pDh#R}�Y�{��%�r�� �.[��M�g W�O��/�:w��)����|m.����� �p�\��q�©_YG�.�P����@0�������,��eotCf���,�£W{�ɌÐo \��,�!��t�+v�xV��ud٠v���`k��M0�ə���gl���u����E2\֩ɵ��Z��N�X� �[u6ɥ��ܨWi��@���8BG4���b�� �j�dW/��o�7w#=���CڞBD3^�aӜr'N[Ҽ}��<�n�4��*I}K��\A�B�8���������)<��
��� �;�p&�fB�.ĥ�;U�f��3�h=�L��a3q��-ń�/X��B���B���H����T�?(�ߴə�7�F �xj����F��O�՞j���,m�mn����|�v�=!��������{�˲��
�LX����wod��l����n�'��i���C�ۏ��s9΋q�B��,#�|h":[L�׹@ms�u��λ01�v�7�;R Kیq�~l��e��IWU�A��g,1�=g�S�0��X�*J�3 �����R<nې�/����h��Aݱ� ��.%�VI&(��!�(nU��r*rW��@��*�������w�	���_�M��]m2�cz�g���h��{���݊��3Oy�=%	���Tt�h�����K��§��է,#4.�T)��K�(0"��z���|��0��6Nm
^��ݦ">(Jn����@��4�狯i�'�E��a4�2�I�X>��;g�
����#���òM��1��4^�*��+��j�Rhpݯ��~K���MhVX`�8q?��x��+��P�č?
��/)��B|m�Թ��Òp�ﲄ��y��_]U���C8��lB�*^'U��:���<�i�Fs�F�<��i�X���Y�HnP��+-��ݾ��f ���|ˁ���ޓ�I¾=�����*&�xO����b��+�9+At@��!G�����lo���|!���H_'�S�����5�ǳ�ӑ@*p��\U2�jە��:_�������ie`F�9�L����j�+<�S�^C���~nJv5�Z0�}i*��R�;b���6�����Զ�c�	^'��d� 
wRBE�V!Q?�i��y��ʡM�\U"n�lj�%����Ww����+d��'�U1��|���q�u�8!�O}����OV��9^�`a|���4S�v�R�_Z�rX��$@�$�Ō\�{��?�\I-�_$�~��:�D����߸�,����q���|]h���V��Q�)��|�_9 $�|l*�����v����@W�罨`�%l�8g&Z��J�	�i}.𙲢xϪ6�����b
4��t櫋���avڸ�v|o�L�: �� ��ʬ8Ѽh���^��8�$���#J��l�Ȥ3}���� �o��I���J�^���ʻ�}�i���Z�[�(�y��*E�<uǚ9#�75h��%�5'�=7w h��4���u�%1���*���3R�o���q�K3ae��{dn$x��뮹�ܥE��X�ľ:���旳��zp@��,�k��9AJ�� D?�q�;��W�ۙ%M� J�0r���J��'������vɤ7�	5�si�#e�a|�;�m��F� 'r֟���ӻh������~N���Mv��,��@�Aeא�0x
���$��9�W�1��8�z$�%�:�&�U ]d������p/�1iq�>�wʌ��v_����|D0E{��h�_�{�X�~K�.*dF�S�hB�k��#�ԩ6O �A1,~Y�C��t�l+^��NΊh���j�2��8�!��x�N�A���ee�I�x�6Z�R�3ģ����Z��F�'�����2��T#��4�[�L1y����L]c|c�Vҕї��w���
��$F �y�!F{@$���ƭ���rG��}5��M�C���3�z�^�υ:8�iɔ�OH���T���p��@C�z��
O�[F�@���
ėј��� 05��.��"�t��Ʌ��gB�ӈ�R<;�(e[�������ݣ~����c�=j��z�x�*y��/�����7�Y�����Ĝз�Z�����6��_�~uw��n��y�]�b� �m���p�պL��<�W+�� ⑦��!�L`��Y���aw�(J������s�3c� �!P�u6^^4iY�>�;���T�pΨ��n�{P*�+�ha���Wf�����K[�
:�C?mo��]�Kg�;,�#�	��v������p���L^;���ə�L ��ܚb�N�R��`��=z-�<��-Լ~�G�
�f�SYu�h9����m����ky��3��gH�~I\g�0¥-��&V[�F��49�/��3d���#�A���􍨛�\��T^[�ђf�^-W�g<�%�
���Sjp����el�Q+��pC~�}M+t���\���3�|	>�)��]�~�6�����Nz��P.Fc�6��W�A~�q�p�����)^�d16�/���� ʇ�u9�˭��Ɯ1�t�7��D&d8 ��k�g>�9e��h�����nwX��=U��������ӑ���^�n���z#�?�gK�Y݀\wd!�)M<.�Aj�_3Nߓ��s�~�"Sj�Wt�6Vm��g����-�J8x�d���U��Y�/���	�� �$�G�U��^�z�eA.,�7TNF�6q�|�h�48���E(���2�]�h�a|��IK��՞i9T�+d�TZ������Z����M'}�f��Ft��J�E0�W�x���t�����T��
u���z��l��Ct���9��#��/e���3k9���{����W�r	]�vZB�R%�i��Q�!�q=J&k��i'��|��#��:�5��B	�.�(S�9����\T1���Ǖ4�^�����tö�Pb�An'�p.��2�>���b:К��-}��P�x�zܙ���~�Z�0�D���[�*�z�C��t��`a�����S�Q�C������$MBP��v?���c�ΗSBB��WC�ol����4�u�����0�����,����:�n
���/c�>��#��������~n�F{"	�M��0�J�ڋ��Y�����9L{ٌ[x{k��)қ�P�nE@��� �@�^	t��c#��ڣ���*;g~�/g��_����c�r�ӝK�26	�3�kOrM�I�c�k���b餍,{5h9�m��X0AU��l�1X֜f%p0��J��[���{U�SLQ��P6��M(��#"=��U�����X*I]�]�g|�8�c�V��
6fCC˖��䓂!�� C�4�rZ���\PBE�&�d�d�n:Ӣ���%t���<�OG� 	�ͰX�Nt�hX�#�g�ݣB+nTw�V\�ݽզ��`��)�^�]$@.ë��M]�s�.�ԀI�\�MfD[��7����?�2' ��0�/����l���"&F�H?޵fc	����L���"q{�Ns=�e��{�j�0�~���Y[��c�6�R�) ��Ʈ�c�Ɣ�8�6��i�y[�!�K�v�2��������|1کt_�$�Z�B����