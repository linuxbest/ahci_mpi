XlxV64EB    26e2     ba0$�ʖ���Z����>���O�Lu �)�L7K��x.2��*I�b�_._H,_h�cL��3{0�:d�7���Tu6ݸc��@L۽a	����3S���yDw_�[�~[k�[i~1�_T�K�/�-����0��5��pe���"�
�`�akR�g7w�*xS�s #+����C�up���]&�H�*:�;;K4s?�6SƷc���n�����I?�|�_����v�+DǬ/L��<����� �u\�GM_D�o�� ������6a�Ƕ��u)��qkM7J��G
)**s����3��x3�},r19�X:�ݼ1K�2�L�����H��Jt���4�1��� ��+�s���jJf�.@Z}J 2��d�5P��;�C.)��mg���ɷ�.pҊ:΢D�H�H^�:ۑ�6y���7�����tW����� �4�W����`R6���{����'�M�:c,~�����8�xw�Z���� �O\>G���2�*�I�d�R��	p��+@3UEd)���	�]~��\����$��pvEny��M@w��#�6h;�u��9֔=2ӊ���6~��G��!��8�쓄�z>X��O�V�4�"s~Weͨ����iD2j6ʟ��k4��-s��Xl����i4�u�C����y@D��pR�H��i�xq,$�~��zM���#�Pד�L�E��hξN]�)��/�_��^:{�"X�X�Dr���Bv높�r��-ۆ��91�,�2ɕ!Vbo�twy�!� y���/B���ğ��� ��q�xҥ
>_)��Ls�0T*N��3i�~�+7�	�$r�xb�����O  ��.��y����@n�[������3�<2�Ӡf�lj�QT�M��(}�=""�ޞj�D�W��#>C]�xr'�����9�a�B�{2�Π�b�8ݑA��lv�o�2VPJ1	�ԃ�P+��mޠ��Z�I���o0��j����{cZO��O����CMd��M�<��J/�nлА8�+�~�2AJ��4��M|����G��$6N;gÝ�-y!�*���+�/�H� /���]��m,�C�T�Ǵj����`AJ�O���8�:yṴ�٬�I[�2�7���LL��_�rvD[��rO��%���1D��`�&`bV��I�$��׾n�2�S�&h�[ԝoW��m�0��	�O���!��`�� �ZE�R����A���g�{�h3�'���ԣ�^'i��szn$w�7v�#O�l�]��.�[�����2S�9�>2W���%x��,�P��S����  �ʗ�ƛQ��$7_��] D�@�(8��N��t�5S�b3��D��[�,#Z�����˟\���$o��^��By ��/�}��$������]��3�t�M�5F�)�ה�t�-���$s���U/���$m�9�����Gaܛ��W�b�k�*�^��y�W~��[�B'�K�+F�����]��a���ouxX ����n��H�p��EAW�|���0En��O��r-��)P�-���oq��u�
�TVpC���E�|v;�W�;�4Mۮ��_41ќ?Z?�n
�hsg*��a�6�ذxi{<����B˲�I3���Jb_0�g�說`�
�����+Kqc!G�E:VwS��V��"c19���+�����BȺJ�)�^��B����xS�K,a�Qg�3���1���,�����Q�,=Aȟ��FߑM��O$��#��M�}7 Z��5�� ���P��@&�C�g���qG0x�w��f*�Պ�����lqC8%4��2 �,JY]@�Y�0�[.������W�gDoS�~mp��7���G� ݵs�2Ҹݢ�b��.���H: ���/�QT)$�D)R5]%�	��]�ț��$U�P�Cߝ
I]{�d_�&S����l�*�3p�PN@I�J��cb9+�r��V�l�π�;n?Ȧ�ph�`��Z~+��e����Jvpm#�� D����@7i�l�-2ծ�#}l+�9����&�/ c����Q 洵�q��Z��\����s�+��_I��݂\��.�*ee#�����B�"y����`Z���b�lM3��c�#�ac 4{#��P��<�j����Z����K�U[��CL��Q��_ީ��d�!��FVd:���ɿ�鬼X��m����9.�8�q�yT��:�w?��>wl8�N��68 ��q��\�I����y�;&�^�Ϗri�ܿ��}U䀘�KQ�<��wB���f��8�W�\�PB���=��Q��$;�����''"�L�r�ݢ꠳r�ú�瓕���\�����p�U���ÿ�o�j#��e�h�ڭo�Y�,��5�Ԝ��_E��֞��MC��>+�y�!���f�K�:��B��<w�P�y��hkg٫A��cB�̶rzV{���#�����c�V4���}R�6K��ߍ��$�����h�����yG"t:�8������}[9- ?۴`F��u>�x ��!�:��GП�K���(f�z��w�Ƃ�^�h�B��8��B�B�5�q)�	��BoF�R�Xv߰KX�FV ԕ����8�JRk
ػQ*_���B,����AI��9�V���#�L��L6�uJ�6d�'�@n��b�Gm#8ڄ=^0�{�9�zf�j#���@!xK��|���D��0������e>]��ua�O��G���y���1��8�*�$��J�T�`Oо>0ov�+�"s�U=��$b����IC�t����U��Y�$6!�96�U��:J�0���&����^ �7)	�%�k�k����9X{�uAAy���㶠l��A"h��=j،|���0���m1��lY��QC��~�,c��fND"�&�E�7Ld{�6��i��������_��|�,�*��t��0M1�ڔݡ���n���I�Ԕ�S+I��R