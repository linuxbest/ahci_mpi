XlxV64EB    5ac1    1280 `��t*�/�OȤЕ��Oq�0�췊�
�UD�	u:�Bh�������섻�Ҙ�Td�X��3"��)�9�lTQ�7R���s*o1嚻����k��'�<�X�t�xG1���N�R�̭��g;�^��
\ƿp��&��!��_��P}.��ׁh��q�$�S̠.qH����%b�7}�\h8��y�����=}q{`�8ʢ]	٤sC|[�T���ZA
��2�(A,���v�T<�x�8�6�������Lb�}\���ww)��(
K_�����8N��h,�5��cX�FЗ�h�1L0�u��o���|��&(9�W��
�o�������>���\?�������(�a�]ao���k���T^Q/��'1��YIݰ�.\��[�wV!!��w����f�K�����"n�t6B'	�b�s�T�B5��8M�%�G<�Z>� �w"i�vrt��"��ڳ�ۮx��]�J�!�����a0
���������;����h��jk�,W�����>��F'RXr���>;��,�5�����i�t{n��׬�ˢ��3Ӿ^Q|k�|Uؚ���{r���e�?��d�)Pb4y�&�,?���'*���!�X#S��vcP%����aw�~�wU�`���Rq�0�|3�K���*����Pl�����=�RQ�8��^�E��T�����CH�0�y,3$���0�4����3	�)���f�a�%��Wa����<��8[��dÓ�:J�CG�U���s�)�;�riW�4��7��'mI|^}���9�t��>��d�Ҍ�ҋa�����ф���v�=D	�Y�mM��+��QT
���z���v�a���H�m�5������Y�N�5���Mwa���;��G��z-W��O %�x�����-9���	�m�R����]YC��b��}t737	U���dS<	p%Պ �C!sgYО�n�T&r�BQ���tS��{�d��<dKG�� `�e<��e���S�B{�X�_ mW��z_�^3�'��Y��r��Te�Q�T>����s�	;��23"�f��]^_�ת���Ha��*e�i�S)�4�l^Kk7�*�;A5f������K��PƲX&�-ՠޓ5ew�^��Q�ðv)���a��m5��C���cɦ=t�	�X���-���|��ϟ���V"�n\�>�b4e/Gŷ��r�+n-��Z0�+�n
�g=����~�L��	�%gyNX�x=�+�3��48۴_�?��E�7�}+��'8�̽����
8�VR��զ���Pm��38�����(k@�a)�y�(/����'�����3qZTL;#	c{����K�D�[���07H��bZ�]��<|*&�Zl�;�9eL�j�V�^��%�^�W��k:���at&[�V�oR�"a8������KCޢ%1�FtsF�ڲ�8��V<�.k��ag��kbˑ��%7v�k��*�k�PYB�s����u���OɁ:�3�-��%��4i�=l�rxj���1��V�{��x��2&q�|��rK����_�`�G�h-�Dg;�5��7��*�Y�[�/��F �aWU�5�g�v�� 77N�Β0��`��r�;�<��]�q���������	_�	��ؓ����<��\���ִ=��j:@)�Z�jS5�^�y��^ٚ]�%nڳG9"&��������l~-k�1SPA���1��@e.���M�Y�w���~���c�kZ�z2�T]�׬���_-Y�.��m ���P�7�ˏv�R��O����S��m�����V�`j��t�|o|�8�d�ruL������G
-g8��Q��2��,H
q�?����4��'��cbrI]q(��s��zf�t�m�`�]���SQSV�y��=#�RR���_�׸�v44+G������PTFxM#ȭ��H�*����\��"�u��f���f�#�q�;`��+�������6�,/�@W�AК{�a}i����(kw�*1D�yD�1::�"$s5�+\Q�0n7�����K�c��R@�g}�¹dUQ��R�?���ź�֞y���%��)9�Uͳ'/�Σ��o��VpEo����Ru#����Ȭ��s =����`�N&N3A��3�0���n.��0FľRP�_EHi�Q���u�*�he�
q�BLCd��E�e��_z?������w#ǀ�sR��Z����uF��W�P��lM���V3���\[hsT�|���g��F��*{��?�8zn���w��_x����˔s	��������&1|�Z�لkT���	+�j��NP�B.2������}.`OXz7�`�x��\Eq��{�z���+�T�%u����M��"<Se���OԨ���+.��$@ ^���yzj��3�j��(����(v�8���x:���$Q��N�������(�{��.R
���i���y����a	�ZD�Y�=Y���^q0ʗ���#� u�pPl�&T��#۱����N
���k�8��W�dT�r~�go�#�g�
Ȉ��y�]萛�X�y�f�_�����)rD{��Qў&u�nf"�8���55�ʈ^}DU]��y��I�_	�j�Ys�Ԩ,YAs5�� lʁL���lF�$#�R �}ziA�Y�֏��~}P�n��BF���0�<���kЧ��a�y��|�؅�%�b"�
~T$}��Fj��STd�/��'��r|��1�s����T (�ԦG�z��cӝ��QimجmE�����9�g�,~vb�5��hEÌ���dKN��(H���9�:����o�y��+�n�)^�� ��Q��T��\b��<��ޚ�g�mF N/�U(U���0�|���E	�5�h�^�8��;I��1�LXP�c�1���Nt�W��ٜ�+#KJ�ܠt���W\vG�U/�w y��"�	P/���8SG�1�%�;	A�aw�����������CD�F�7H)�,�Z�C�*=�cG�����Wc7���E�9J�[h8�i� ���g&�ѣ�Be��	��ʵ�/���5 k���Q�Ha�W�w|ׂ���5���9
l���܃�
��ˢz`MC�#gTB����}�(��sV;�.��`��n)�'��K�F�*<�B�`�{�zh�#�e�7*�㸿*+�Bª���ܥO��ނIF���HKp���}�]�r��Tk݌q ;��A����;�-��<&��.Xw$����t�P� b����U�Ӟ�ܩ��bM;1����a�o�+Q#X���3Kjr��͜fޙ�SД�<��� ��/�}���M��˯�L��tj�YɝY�(s�ʪ٤HTx.�e*�!nf�~�d��aW�����j/7�|B��c������ �jݢ䏼C�_���WG�o��w6�>BI�/A�P��9ƒ���=_uW*����/�D�C���,!�~���,&��/Qg����k�_�:�-pj3y�Ƈ��Kcn���&��?ب	�KyX��$G��=�J$ƭ�;|f��6)(M� �z�G,�Ƹ?P�&۟����
�@��P�O��Օ̙:_Hъq����9I{�״R_��&�°Gݥ��N��Sy��*���>��4�A�80�DD"�^5#{w�FKd�wP �(2�w�Y��o���w��r3��_dSy@��C�W�\��;���T�����9w�8oy1�eS=���!oԂ��ȗ�j��1����DI?�%���2��je�-�c�.�ɭ�[ y���5�p�#�n���a?dk��߅����O��џ"'�'��
Q20����!׎��#��l�(_��p�*�:u�w���2xd������Ht&|�.�n�����['G(D���`H��O����;�1���z��zJ��T�[LF�,�	n��i�鑊��Ȓ��O}�(7r��G�A)!ܷ�}
�&d� G�n#��7xF���K��lOɼB�F/�ͩB�(2��5�J��Wy�"\���Y/��3̄����~)�|7�����^�f��퉛��G_nS� �Ōu���!��S�f0���M�;� .�ȤV������y�7����{����u�������Z�T��O��A(sQg���B�n�D+m�W�6�J�d,��W9����k�6C~��W�W�Ղ��-d{�e�J��6��~�ʓ:j(� ){���u��������͞�6?��`x�}�C�
�=���_�F��Ja�	��@Z��ԩ�0zS�����S�)������MI!#bH;Y��h|a�!fEV�'q?	Z/��B51:��4�zG���~�/��Rh%�_T��q�$C!����&�?ٹ�J+�H�����vR�H�Î�b%�XS��KU�7V�t�DM���� >��B���;���YX��Mƒ&��!���N��,�ݜ��n��}�}�b�a�k$v�%bS>D�	�(n����&��]��01.��?�ڛ�R%��L��K�c�NA�M�V��%� Z��?���jI�8T����?��a�
��0���gg�B���$�!�lI��$0j����Ѥx��r3e�s�,+�B)�  ���p9����D�����i
�Ԡ9�X٬L���7�P7�	�%��G�%���� ��o�5��U��N����Ȩ