XlxV64EB    19b5     9b0%����~�n�D�*��\ן�ͻ�+�{�}��}���i(z����`w��S�Z�㵩�'�߬�%@Q����q�b�&Ҥ�z���H���Y<ԓ�ݎŮ�Gʭ#)�#��o�?(A�e��T&���Y��u�i�\)FŊ��rS���IZm_�X}cW[zT��T�?c�S�K,��%������r���^�'�ˠ��ƣ3Ÿ����^Y%�_�Sp�%�����*�^~7�b{�)�A�mբ���_�mP����1�$�Kֲ%���U�V��0�81����pWY�/�>-����H�z�6X�Fk�����O���U�	��zևe��0?�����V�,���d��.�%���N������8BH�.�iRgI��Mk�LF���.��#�m��{�갑*��5��_~��k�$q���f�/$i�(So8/���	�Ч]`���q����7��^��z�7�q��\�Y�w�%m���)��ߗ3��B��Y2� �܎U��1��,��.�jXa��s���>��D���=�7V�4�>y"o8=�Q�3t\r4a �_J�C�Mg��Q�{	�� �ɜ�w����hm�J��
ۘ�$.���X�E-��n�K����5�&�S��O�:	6������&����_��ԅ���o��5ƒ���1����N��?��|��� �I%�.
�w����uN$��i����}���"��GOp�ڛN~6\Y���G��[��Oc��ӑ<�����P���y��V,�N5ղ��U�M3���Mu�zj��*D�{S�g�Wp��c�>�k��f��'S��WqD�8s��<�q��Qr�e��c� o�I�ݬ�Z�4�����	j[�ݏ�A�맃�1�Z�,S�|�#c�����v�C&�b5d��ek��#P��;�������ϝ�n���֐w�=̉�~Z�|�����䩇i�7�wi��^6lp#7�3'~�D��{���@�Rd�Li/�������de�m5�??0U=��n�	AOQ�l]$sc�@n�]�1R��3�V���4�	9�@{[��s��ו��9���(�o-,F^���%�3�2���<�bDiY�d��G�k������I��D��g��C�W�1nU�q_2QO"����H��h'�@��;^����wS���0��y.��!�U��<��U������E����J`��3s��pÒЌ��,�.��@�c�L�����U�I�F�,�8��G���Fu�b���"f!�Ԉ^�-`����}fe�/�
���s�Ԣ�+�����������
?9�?�����%�Z��4"�J�r��@��|�kx��{*���q��(;�����BM����������f��7��e����:�h���FP�S�YX��p�@b��X7ŪArs��{T�Ӯ��w�շr�d.����f)��;je�`N�Hr�-�Q7�*ő�GKn}�U߁~��K��#�Ȳ9섹�hs�����`� ���q�v��r��Z����"ax3&�_��a�z�I�tY����]?���� �P�*A���태V�ƿ[0�4@*�H�J.�i�� 2��:�$�Q�o��A��g�LI�`a��N�I���p�{%�7F�_��kF+�j����'����G4"�*v�<f"�${ѯ(��}d�{�Ɉ}��g;��	1X���-�"�����?��Fu��'�4������i=ٛq�ʐ�x�����J�]k�P�S�_}e�y�rEnܵI�Jx�mv����ZtZZėp����搻��+�qe��5��Y	7���D��r��K����9p��.�o�_�ᱼ�TY�9V�:]�~2�F+=�H��=)���v�#%&*�f1Wj��N�+�KT��I��;pv�|���&v�r//I����P#X����M�/��'f	�����*A�)���ԇ]*y��kˮۍ����v�_3G�P�Ey?g�n�IYч¤��2ITc$�Ib��dO�U�W�a����h��ƍ����bG�UJ~�C���ޔ�@󤰂ݶ�i���^M�;�����6W�ct��i�g�U��/v����B��kk�"�N_	mU�H A���%���P�����˂o���.��O�?��33Y@��X�qv�|������1/�J�5� ���̱_:}�@Fwt��\t�[�r��*Ư��%��@+2ӳ�����`x�]�T{��I��Iencrf��\�׾� �Mj�v�CU������A�#�X��i8����ܦ'Ee�n�6�h��L�i��P1��}����*K4� �,u$d-}�YB�M9Cr~���Y�w(39���!��R ��G��� \�:��Z��K��/�I��-h�d���i�'o�lEP�Xd��{]nV�^��'�����tx]GV#����ά4��S������I���e�%���