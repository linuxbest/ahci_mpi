XlxV64EB    17e2     9b0���&QA��y9{F�b�����4=\f�7�E��ﰇ��Ґ��^i��U�\�r�%����f���/�PZ����{�L����J���Y���� �qO�~�GV�z���4"�o�o)�Twg%(ߙ�c���R3��ٶ�qz��9�[Hu��'���vX(KݘV���p�4.�����4��UԈꪂ� I���XE};��|�Խ��[��nso`W�ź���S�EP��;e)�%x�rװ����)�EI#�s�%.aa�����=�ڴF����S�X;d�VW�=
��ۣ�A��	��۔�����E�����$���a��2C)B^��_��7���M�7�v�6�a���)���95����q��%A��M7��}�|�'²~1�����k|�+1�p@��J���S�ɲ������Nk+�3l�U��ߒ��LuU=,8�a��/o�I�V��2�>w��i��*,8�t�};��i'<�%W����9� /cN�r��� �ɹ�Q3�J�e �*X�����8�O�'�x��o�)w�CUm����S�ASܽ��^��¦��ϥ�u��S`�T Q:���u��s�XJ9��Ҁ�x-#�r�fA}�f����+�	!I�{C�E�\��r6�0f�a�ؔ{�[Z%+9Np }Dh��"�n�?�`�ݧ��K����a�!e]�4&3yƄ��W&#}2��M�8�o���g-���f�Z����WW�Y/�*̵��T�'#���\,�BB���D�v82���� aM�;�="�E�"I�b��~��(���,����%��z���=N���Q���>ٝ��2ek���I�&����]SZ�N ���"�^�92�=��͐�?Xa�\���~�9���t^�t�-��wڀIQ�_�˗ޗ���E]��(��̴��j�~�8�� ��^�Ւ���ld˿|��l�LX�r��f���lT9)�i׏�.�@��K:��[<��noX9bI�w�� ����Iv¹oz���NG��X��n�t��MY��� /��뉶����9�93tU&&1��L���x�^qtH��
yF��~>F��ʊ-"L�x(Cܭ��0�
-�QW�Y��g��Ѥ'�\&�Â؈��-�ޒ��̮A!��a:�A'���>k�<_$��'�A  ��gG� �k��ٕ�;H|�P4$_�xS�3�D~<ZٷF�3�q�V���SčN��x�����::MlF��4t�m��*���UU^��p{��y��_�
�M�,���k���$~K�������2��U�H���JN4�Ǧ��@� )��H�m���= K����8s��R���7-��Z��ŷȆ�����l���~p1�P�z��|���Ze>|��P��$D�,C�)�ߒ�Y��j�y�+8��AM�pk����9��c����KP�{���˄yF�{���E�Ű��gSi`��y�I�ܥ��e�ˍ��~V�2Q��$�����½3tI�	�ғ���<��; �=X��/i=L��$�<�.��?n��@0�Hc`�����xb��s�+v�ދ�ӪCþs��2ӝ?S�jX̊��9�~h9�9�i���f�0���w�4ּ)$�w��0��髢�d�_pa;�h]�[.�� ������4���h���M.���Gc*�X�>$-Ͳ8
o�+R��у���/� d������i�1۴�c���N�Ci�ֹrâ"JH���rvh�k�j�" -U�Bڛ�[�i3�����-�����?zC��9.֞G�J%̲�P�̲G���
��5�]�*x�ZB=��Y�a7��a��/y-�|�8�)!`�b��f�Q��[l(�W��pkB*�P��KJda�����+6l��Eҟ�E��K
������1+�fM=��D��A���:ki#�rMT��o�<9�� �t4 �T�e�_���Nx�YR��a~R�G|�)R})Y��Ӹ�Ag� C���B��U6�K�I��O����l��l�<Q���Re����i#�giC��þ�F愬h͞��z��o*��qJ��Fe>U?
��O��[]�ZaY�E�r����r���'�K~ �"��t��p���8��f^�z(��v~�T�N.aSm���������!N�f� A��	���r���~}�ۂ���:�Tܙ�sЗF���Z�>ioq4b;�%���Y?/@Y�h�k~ #����h1'���Ц�|�٨z/����k\{yxV�,	:O0�4G"y�~{�%�S��Z�{Q^�B�f�Q���W"���@<�TO.ޱ��h��L�m��b�5Q��Kî�t�����KlF�ݔ�����#wN�;�"B�}�!d= �
qFIje���$�9����g�Ŗ~�/�[��8#�(�����N,KzU�'����֍�9�?DW��&EP���%��y(߼