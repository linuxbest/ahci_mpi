XlxV64EB    55c9    13b0+��=4t
J�c>��2�����SF�ʔ���d��l`�o�
,?��d{�i;2&��ϳ�4��:!��%��Z�ۙ���,~5��S��^]��� 6[����b��[�ށx��)[�O�k�Ȟ7�/�,��iAѫt!Z�}Q\��ËDѤ��J��YB�i��"��$("��&D߈��"�O.��Nb��`Ϥ�W`��Z����az82W�!���9�� �$2�(�^�1�<Եst��c(�f�h�a��"Ix�e�� g6/�s`��[�|y=
Ow���%��"�z0>���(�N�����\��m�x��3D�{�y�K����T�������d�K�����z"E�Ю��yk
�P���K�jJ>����<��۷\f�J<�'�2j�lF�}R�k,"z,j�g�)��U��N�ZB�~]c����q��\A���K|9,}P�;kKі%Ҹ����%%w�����>�7oS'dX��5/��xW�3/Ecո��۪�v����H+�ju��B���[���
��0 s�x��������6�?��ܠ���ʐ�c,��'���/PX�{�����B����>q�N�{�?�d����=�z����n�L!��`j��*z�˼lb��:u'��T�\�~~�}�A�ڞ��h�Ղ^/R�m������J�V�l�|��A�3)q90��疥cz~]v��<ڭ�gS|��w]>G)
=3���C����B�	W�~U+1Q���h2��*<�}*�3A�!yS�ƌ��O�>�N$r�t��'T���������P7�*�!�b����� m�:$���H�h��'	��oѻ��2�}�S>�Iޅ�{z`wW~�3J64AJ�ň7vW�w����RoO-�%AIƷ��O-�
K���A�6���$��N��xL�r��m��[�?���ܢ�h�.8��	7Qٌ�<���iЏj12�ÂM���|��Xa��#��N�ﳻ��d�"�Y��gt����/����А�z�N}5�gi�Pe-e���d\��4���)���у���;鄙ce���X��'U��]o���E㧪���B|<(3�`_��=���������������qE������A돈�k��5T�^��;��H"��Œ�e���(��~��F*�	��Js`���b�}��,������J��-�<Q3��W�$7!�A+��Vé>ZܸК>�{:�(j�����%Ҵ6ݿ�;zڊ�P[�
&����*u˘�}�C� ���Z�;�%o�F����(K���O�	�Hm.�fB�˕XH���(=y1)�����R/+Ҁ&�7H�^�o
b����!�3�v-�~4��G���jM%_i�������1���+ϔc
iyV�1��c�qn�S���D:�P%�*��^4}�/�̀��@*m��a,�A��<$߷�-c�WN��J9���d��_��L22#��$R�4��s��m�7|�4��<�u\���qb���(�I��a~�Ց�Q�`x[�"�?V� @����E?I�i����v̻��{94O�/�F}��n�daXZ��A�PY�-���Y�B�}X%���fMJj�ψ�X�=a� Q�h7��H��-�Za_KZ��]�eT�a�6��+�S	�:�K��f�(���X�s/b�,�K-V��^���n��q�/6�A����l|��'��5!3l����ۼ�;��o�LF\2����M� -���� Q�+��q��&u��G@oD͋��&z�
�I8�~/��w�*\RSx99�u��Z�&�?�˳�Oվ'��9���o� "�0����c��0t�����n�D�(c��R��~\l����2ڂ$�/�"!t�)�:�C���m{�I~��ˆy%'ӓ�t�{�c��AZ�R�٤q��?���,� ����a	���t�l3N>��5�;*>��zZ4�	�-)�>F�fɢ���5p��SV���m����@X�_���Y$�.Ī��I�2*��ʖHeR8���Sm�Ik)�*x���2Oފ��_��mӼ�At҅w�\�#ª"����Σ?���,55�s�ۺiK�-W����\�@w�������5�����jT�y��|"�X���֣�-t�t(�:��x�*����
�ͩ�=�i����C�tȶF�-ȶ*S2�	������E��ܸ=�"gJD�]���^HЛ5%�žT!�'���@�����՗���M�;$y��;ʕ'�UF�՗�6gY��I����0���'���-��H-�(��� L��vյ�@J��9�,��rD�B��%���B�����4$Q���>F�ޓ͑��ZN����s7�>���۽�Z7��8��'`C��gx~3��g�<�N�i����-����z�|FEY��(���$D�A���gQA���4sv^C��Ě�o@�fV�_<z������^U�+���Z>��t��E?���w;�E}�|բ�Aa�X�"͘E�����"�A �0'	����o��X�F��m��e���������UbZGN��M�j-�	�}�����n#�C���=vR���;�g�"2�Sx�1s�@��@��}��Pwg̀�7R����6�'O��P��.�9�pR�`��wi�����c�s�_��&�U���/8�ތt��	���qO;C%�=�0���?�Qn E\kx~�?@bJ<V��\�s�f��KڬG5���	�~��A/s�Hm��p�#=E���T��_�S ���P��ݛ����V"�L���A�j?��U�)B�l�oT���cq��g:��Խ�D�@#��F*L�hay��T��"C���m�ofz�Y=e��Z�a:R��6��BQ^T��JzyD�)m��_b>����[Ft%����u˿lP��T�^���T
����pA.�٤q�vr��$IF���/�q��MR�ᄤ��arP�[��^;�G@�#^��36 ���#V����(m� ����>�� (?QJ[�l���y��)��e�j�'9ߨa��m��2`5�$HV��d��P�DN�RV0���s�!�4$
E�hY $�H��.�h�$�ZU�:A�ݿG`T��,�-���I���d!I�f޾��2�$~&����kW ɉh9M���o|>[5O�A.��F��>�O�<�D�(T�K~?af�c!Hl��Ⅾו��X�V�^$��6pwS�G9��b�>��sU�VJ�@��s���̒���Ƌ� '����8o�	g�?��ř�2]h�m�o�B�����h�o�"T�}\d{M�=#��N��XA�N(�r'����� �L�5������Kq�P'&X"L�hu�e���y�n�ĵ��|�V����R�#!�?�)�@����!��ŬfK���'�c����+^0���i����ڽ\�7�e��6����0Y��$d�^��ys�ס9�Bڝ����P�D�B�'���2����<p/�C(6�'�� �J6���X�EaG^#&�9�1��kū5 ���cs������ޯZ����=~���Q�Ћ�����|Η���3����G��.�t<�8����:���\�,�K3gU��@~����5?���(߽��TiɄ��k&�\C����gP��ҩ�r0B�m,�w��(� W�*5��b~k悚鿻��U˽q�|�I�О��c���@���4s�?:\��Z��:+U�?���
�ÈK�e���W�蟄�r�t��Gt)��҉a�.�dc :��#��}teX-���ӾetϏ��T�n�hp}Iq{���,u�q�ĐI�ׄ����L00�מe921nU�;��

�vq`X搇��:u �<Zb?>����@4��3ǧed<s��y[s�r�y��)_NJJ<`��y;�����Hlp%Ɍ�GM�	��01 ��g��ف�ŧUym�,4��vL[�G�B��x=s�.��ů����U��ٙQ��Jm��k5LnɊU�*�=��Pg��I�Ngi�\��:�`6�A6�b�B
t�S���'��m�C��k���4��X�p�J�����*������|��i0�B7�ppB�4C� 3�����߄�j�m��D�Y�l���P6W~��Fհ����E�ۻ*y�~�'�N	C0,�����{p�|K��?�i�q�H�g]� 1 ܵ<8�	�0��:��O�ݞ����Q�l~U�@�����L�9��q�Z��R��>QAJ�{(�Yl��|3{S މ�	���W����	�T�"m��@��p"�#������絉�$�c]�q��+�N��Z)N��k����K��8���8�^����@��{y�Sr���ؔ�t�Ϙz��#�em ��=����iӮ���xwh���c Cp�J�١���K���c]���!�ڄ�v�s���b�}
+�b����굳�y��[��f��'ȣ�O~	��3��1׵M�b�S�,�:P�̵�4�P�Y� 9���v�O>�i�<�K�1o��{�e�0K�Zڤ����A䆲5��@s���5S͂���yi����<�]�GZ0b�+�&w�359��+PؿDs�9U��9PۂQʘ��<�
[HV�J	Og8��/�'�J���b}7�����ߪ�6`��u2s]�]�U��7iY�v^r}��5ő��>9��/<�(ۃ����X�l��rv��_h;��5�pq�-�C��Fg̒��;!��.��yp�D���՞n�8�}�9`"�y-��;3��t"wo��1�n�M�/�h��sP�'�7�%��kY`��6���i�;'��e�.B�%�'ΰ^����$.B��H��J��k��h3�!Ϝ�B0�-�F>ԩ�qCʶ���Ŋ�$���ߋ�@��W���0J2L`��ֿ��b|8�6_/����:%�ܜ>�J˶���"���U���w`��ܨV�����MR�"��x¡�U���Z��OZ����