XlxV64EB    5891    1450���pX�'(4N'ؐIp��x�A��_�p`<��k������q��ٝ�R=D��k�)��_�^�a8�ڼ��Z��o�௢"z��3��&#ux|�&��T e����!����E��������ƞO(��0�ۉgK�8�A+��]�d�����ɪ�M���x�X�:%��*67���ҫ�6wƜ��BⰀ��[Y����ޝ��.�İen����	�R�1pR�T���/b���+SL�KK�.���Mf�곺^����Mi���km<d*G~%lQ��a�E~���ω���Zm��1�<�ZK\��[�rz6��ɿݛvrq;S3ڻv��xlR��Q��M�""�G>r�BLl�L�W޴�
��z	�㉶ǜT)���(X�Ew���1��4dVb�Sk,��A!��VW@����k�E*
|�%X�΄�����]\���W08b�5H,�y��k>x�*Wu�\3 �%���d��%Dj�+1$��}2��}���	 :e�s_k.��=��7�L[�]xIo��B���r�Dj|;�Ӯ|s�b՞�	��gh�( ��Q�fa��ZS�f�@a�ag��sx��j2�XUw�l9�I��|���ŏr�G���^B��� 4$�Û��y�A<`��YΚ�|�b�q�*�����$,d��	���<�|9ޣ5��'h(F=���g���0y� ��ab>f���z�p�M���� �kY�����o�N��MbB�${�1CsHd�Z(=����X�=���w�`q*���$�:аۊ��63����ys��V��V�ASfϿ�;V�m�\�+f7Ɛ�������N�å�a	������O��L��~�E���a��(R�T�k�����L_�r�)\�)1�zV�,�h�[��Qr�d?מ�����.L����ʳ/7�ov�� ��͉Ɍ�F��*�%&v���V��)�`��.�������N�OZ,�Ŏ0ӽO�����u�� �\��Z��YD��9�a̒9�ǳN<R ����M[�u"5O���%��+�>����u��?n �������-Y��~�$�h@/�g�(��T��g�ן���u��f2��D�st������җW��5�Xl_t�!�.na�xhP��	%)�����iu�
>�v���r�iŋI�;w~أ�F�	f���i	-܎�ڇYc&�E�.N:N�!�� �@���dA^�[EB������\[��H�|1�Y���A��͂RB�|*q��tݰ#��qL���h
��	��E/��&+�s��ą	��+F�#ۯ�;���co=��k�m�"��"``n���y�'�.|�,z0(��!A�kO��ml.HZo���������`�*Bc�˻X��bT��	i[P؃�����Z��Rɚ�F��
���$zr�΁�v��Ɛ�%�`ց��,�w�?��f�>�xc����,q&>{�w,�����V�^=��:m�W�D���t���.	�	�I_�}��@]�u�t���_'-ԩ�Y��o�1G�b���O�e/�q���us�����'�N�b�	ո������,r�b��Ѫ�RL�Ł]��ڑ����d�iZ��q|��?R�H�B]�(2���t��=�k����� �����qq	'ժ����h�S|�1�g�_"B�x�Z�Fd{84�3C�Ԋ��\jt!5�]�:�'��	��d���a1J��|��Ӳ��XsL��D�֙�0>n�_@|��Y�:>�|
q�;
6��{ 7ƒw�2�6I�� 
"tv�DY��5 \��� _�[|�)�(]�8��Ǳn7	gY�aT���!(<npb���
���>�v��t/��v���?�7mYQ�{��4aH��ۢ�����=��ܷk%�Ʉ�MO��j\��!��"�ER�VĊIG����T��;�'�[��̖JP"��nʇ�J�� ZCYG/&Ā��iP ��T������[�7���GmV��v��E��L,���ս7�سwW��WqO��^<�(9km͇����_;xl������,��ײ�Bh;�z���KY���h��ܜӻ()�r�b���,= ���.����� *ޤ� �S7$}�>�)��V�D���7���>\Z�*���C��*F���k���X�$?����i`��2���r�~q�M.��;�1EW��īn\br�����ț�ge?*��1�~�.��kM��\O<��5��Xv�׹�lc�J1�Ҟ)c��'Z��������P��Oc	Tx�Jbך"�>�}��l!J�5�]�r��������ch�fޣ��]��C�ҫif��Z�/�/�q�
[ǀ9���kA�E���䓬m�q	b�(�)�P^�׏���7Z��0���[���X����Ԯ�F��r ~
>s�PB@���*IK�O�6� �T'�"�"lL�]l.G�)��O:�I�-(���)���c��Q:���`̩n��y�S.,��e$��W�}|a�T��G�J��%�FH��/�ŕ�P����hܝKȉp��}�q��g�݃nM��@�K��m�⯙��i�?ݓ������Ha[<�V���s��X{��r��r��ӱ�G-=��|U̝]�
�σoǇ.�A&;��yc���bڔ߉�1�*� ֜^{��j���{i�1ײ��PUT��Rh��3�|n+@��%��"d�ԟ�6��dx� s�7�[��W���q�J�&m@�s�J��2?A�F�r���d3H-ʓ_�7��?u5�Q��;(r��;�`s=v�W�C���NA?���K�����e�v%�XF�`�1����.�Z���)C�=x��f��_&�4��B�Q&w���H��F���/~F�h@�[����4���\EϨ�X�"N�Ь���������]�O����xR����q�2����pf�n̻z�T�r�,��?�+GG7�����"R)s�LF����?��'�.���x'=�S<t�Tz֭���hl�{��{�n�ͱ?�CsO�#���Ma�I̙��&N��.�6{���pP$�~���8*�,����u�y�	�W����n�${��ܦ���E�����*�P.�'��aC����"5p+Ҟ�Sܖb��!Z���Ս�K��P�ک�
^����.�
b���׏[6K����+w�b��/���TX�TP� P�Vu|��R�v���<̖ }(-鸳������){�
���s��R����)�1��ɮc��T<��6�N v���Ow����slL��LU���6��k ����wn}���7� ��XOM �2�'�����y}�d�"&�a�%.c�G�bQ0Y�����})�$'�V�E �ޫH�'���N��C~���S�տ��T�T�{g���#f4$��[�Mgɜc�����v��u�u+ #!�s�]�p���H�A��!���Ѕg�<nZ�?��)�θ�.��ԛ|�q���k��|`e��g���|@���f��($��!���%��q��B[�\1�ˊ%9@�!�3�ͬ��V��t!S�g,BB� �D.�H�YA��ǜ���Գ�m�g9SR�.�B���/h0��+���&��uX5������t�yL�z���]�y�GS�� �tc����Q�n��t�M������4H�Pahw0LB��B�����Vw�ҧ�e+�V���@?���d��rЌ���an�YG�Իm�W��d���2�h��G�����)2}�A����	���u���kc��LJ�M> ���	���]nV�g��!�5c��Ń��8}FeMX8����Bztx{�q�[�f5��$�Y�Q7�5GA'������=����d=V�]�u�F� �#"��\<�<Vpt[JfY~*�	�^µbu��f��=�*��*g����K!�K�omW)GF�aK-&�z�­.YM;�S�V��!��Y^&�y�E�*��N[�ÏR�rp�N(0w\��d�erG�w:�<<%V��EDH�q<;_����n��H��A�p�G��^T��L^ ]fV<��}*Q H$�Q�B���6�I�������۷�;Jk�q#YH�{���mDC�iM���1��,�n�e�d�+����Ӧ�,�y5[�HM�˟�L���+��|���=~�@^l��qza�+]n�$S�Q2��ML?'�$&Ԍ�eY��b�R�w/��6� `� n@ց"���B��2J�p\<̼���Hvt�p9�t�U�x����D=���C�mg�(��[�$
 �N���]�\�|�� =]7�/q��w�n��{ST���d&:��qߊX�3+��P��{F�������H�^�m��}�i1��<yQ�.eΟ�X�̆�dg��^Z��8�,�ȕH�4�n"wDmZ&]���?�Fz���A���6�r�{&�D[��}�d>]h9�Ɗ�ֵBZ¢�b-�iJ��x�ﱌ�-�Pa��`�*X��5�ċ��&�K ��L <�,f��_�]��cj3{� ���(5�쾢�T�y$�=m���r5q���_o�+2����8 ��r�4�,�c��� ��TLK�2$~t��6����u�������{���h��K��p�];(#Lk�Ñ�M��[�k�j�NZ�P������H|��r­�dE̱��p
�<���1x�ZA6G��DF��l+<����]޵�L�h�Mѭ>ȓ��"N�V�WR�T)�w!��ow?s����ȡ��3��MyC��D��#��`o���!z/�����XÆk�C��b�����N)_��g�G���[�����j�Sΐ{Z5�9?���^{ #�!�+b�m�s� K�%����r�Kߵ���s%��S|��e�*4�k�G �L���-�Y_�t��M��f/C�����]�!K!����\47J�h��̬f����[a,0��V!�A]�<0s%��+��Km#�%!�ɜ����$u��6H�u���I�I��E��l6a�%0�j{�8�*�J�=��{!�X>:�7�]��6�?_����m����|������)2��~��B���7�D�������٦fm;ạ���
�=>Wq�K��~�ӄ��P{�7�A�YR�p����