XlxV64EB    4a06    10f0XM���-���n��g*�v���}04ufN;,5{�w}�-nk3�+�҈G��O�E��\0��%�a�^ ��OEՄ����bBӴ��2��J1���B�9��';�Zw��@j�1�&_
p�jw��ݒ�Ew�p�۫���u�E���YH��L�����Bg�u16f���?dɀ{�i�����F�����Q;�����r�T�v���`�+�uo�ܾ �ۄ���ѿ�����qaq��վz-��/���'�{��Ӿ"�\r�Y�
�v���돇���v��e7��K{�N;�߁��d2 ?o���c���f4�k3u�V��Rg��wj(N��ݜ��(��(��I�_.�������5)_�/	F�D�CǍ�=��-�9&B��z^�;�̊�y�T��C��wq�j&����9C�a��n��X�%Y�8��o�Je��s�=�)n���E�V��?�2J/ �v�"�dE����������/t�G$>�<ˬ����;�ET��E0����ߢ�ֈw����7�P|4����"6^����K�1�5������S1��u}���Ӯ��L?�X��o��n��e��s�뻟/�dr��~���[L�ulch���7�%�/p%d��L|�3;��<���V�ϑ�ԅ*Ya�~�B��`b� B���lb��S\���$@�X���_�;���"�,8q�&�]�l0zYCݙ,B��[Vl�b!,ǣ��,1:�)�ؙ�w�@��/ޥF(9d��`>q�(��&���J����������E�51	|�n�"��g�$s�c�TLz0-,�|~"��N�c��8��C�h���E�u��H��Xf��l�#�\�S�;����6��m�$7[�V���j����ڀ�]�E��s�)J�%�ȹqq#*ݔ�MO�=��� c�`�Gt���>H��,8�<�b�ȣA�km��6�.�@�I�:5YQ �)��&�;i�p2����x�š�)�3������j�XRк�A�k�l|�N����s����I��O��U�٘4a a%}�ݾ��bu/����z�dX�3���]��~���Wm?VL���9�cB@ae^I9t�4Q�����#�7zz8M�~B��.;�9�JJ�|�@��'J��:ˠteK�?Q�����n�lAt� (���2�>�D��X��)o��bz�s�"t&��0��3g�>>e7�0�c��Ȓߙ��H�ꑝ�)x�l���>�C!(N����D���4[v� �t�MS�:�s`�׆*�0%?�#O�ܔ03�f\.^˭mv��G�N' ��'$��{�}t�,*#����u�5���-u�O�+�qQR�SX<tb��C�h���y����S9�C����w����Xvv��PK*�戋-Y���˯�}�7Gh��j4�\���P���J?��{DX���tL��R���,�D�{�r�<}�%�B8N�?=�~��Զ�:a�Ů
囖P����Ӿ�
�XX�cO�7����.x���u�a����ZN 3��9m�d�B�=?u�ǿ������l�u�'܃T�/F��@!<np�� ��C�.<�ݲ�[�/@&ӵސa8.u`-���;�F��+{�K��P�o�����\8����&hJ�X�I}H��c�(pI�C�����]���ZIX�u���&�^�<WA�(��0��'HNqkњL��g�hvd�?���3�y����/�a5#Äy���U�w���qHa��  �`�������BW��D��Y�<�i���c^l�~FZWbR6���4$7���]k=>+pwXe�_Ұ]J�����}��u��4�f�-�D������_��Q��΀"�5�p�s'�k�UR�
>T��j7焰���"oM��f=5?�4���yq���r�#�c;!�������naYo�̘�����Q��q��.7���r_��=�`�<���.�+$-6�yAX��7�A(X>�^"p����n��b�LM
�5޻bЛ��y~�.��k3�r��x�z��Z���B�M��K�@ak3���q-D�����$Φ��D�*�c������{�d���I3oe��Qx�GM�����U�
�m���:�V7�-k��>�s�h4�r�yMp)����\M�@�����*�)���ٴ�`$f�w�����|�$����j�g�:��;��-ǐJ ���T���j�}���3��9C�H؛H�g4�������,����)l�����`�2�?�R	)�މ�뙋)h����N�T��XUC��g̓>��
hM�sz�w�##�&���8�F�rHh�t2jd@���'��T��H�*�Jda0u��fU��9�/�##3H�����L"�yd�$���y��R��CTf#n~k�Q4���6dym";�,�΅(}��+�z�[UKf`h��(v�Sb����l>iU��`G�o�M��@�{y	HS&��6P7zco���py(a�_��1��d�X��i�����76�r��8�˥K�ۨ,��OcV�֖�V)�T'0���~��;�.,���L���,�E�q��Mρv£ǀrȝ���2���`���f��j�{&P5B�%�o��R�}�t��b�DI���'�����?�r0����ŭG%w���/�e~�I4�՜�=��9S?��;�,4|r���3������V���ܐ~V�&��Ia'��TU]��7 L5���&�pR=�ʎ�U��+��m��?11%�xv�<����Mv.�D|�]U����U�&<lWu�$y:RA24ι��LB�v�ByMi�H�`w}lN^k\�P]!���m���H�J��"��+~�-;X��pŲ�i)DUvJ'v�)�$-j�sA�&.�
0&4쳟m�����#��_:mB*�-=�$��3�K�R�� ��$��4ҋlc���E��l�kގ�s��b5��Emc�#yߥ�\����6ă+B���Y��qq��Za6Mv�#�8���P�_� �A���m����
�|\
>G�}@c�\�?Q�T/�ő�*c�p<���˃�θ`(ݛ�ΐ�~嫭��9{�U�S�j���V�{�򍦞��1��l;Έ�P�h���LW�n�e�P���,J1?%ϵ�M�K�6X�l�+��w�3��"�`dpцQX��i��o��N����;�	�e�J�ړK�O�R�c���p��e�95:�ꠕ7h���tE��mɽy�}8���H-8�֢�f�Z��31���ҥ�|ca��ߋO�_�*_�шn\E�"��2�d���>�$��9����J�<��?�/^�cVӁI] �~�7J��O�Z��P�\s>��݂���(z� �[SƉZr9���nwXn��W���;k:�I�U��2�*������.���Z�@�� x$�N��fN�#������1�H��z������D.�T��9I���\�1x:�c*��[�k���D�ou�+2!��k�d����0�5�OT�i�Kk3]�_d�[!=�����7Z+z���U����~���Ϣf^�E�<.u��8?`Y�lfk�y�5��_]���k�^�;�.,F�~�R��?H_$�[x!��$-�~%)�QP�;(���q���R��V?��c���\_UbT�=]�
X쪒׹�<�f_%5w��ѳu�= W� x�{C�
}���l�U�'+��<{�iO'h�Br�k�N���q�̦r�1�w
��^$�!`Cq�t� �W�ұ��Ґ:���{�M,�H��h}��D��&���߳���3h>�}������KW�bF���C�<��)dL�mF֛=�4��}|�M*8W�A��|����j�&&��^��p����(l==8?u����m���Hu�Aյ���o�5�51 $�b5t��"�&юl�)m[a���3�o=���Ӷ"��VB�>�H�) ���{�������fmA{��11�^�7�<��p<�xɴ�aǪ�q9�pbR�(I�u!h�Z�d�P��1)'�b�Pz�_�M��nc�7�?<>ӎV�R���7wG�V��hn����Z��}�w�׮��T�U�c.���Dh��+q�ͷ^����i4�(��T��u�"����k�����k1���yF�;��n U�ji�A�[����4B�fi@r����gI�������}g�����ѩ����@���1;5�e#�.��\���� K�Ɵ8@0�惌�);բ�W������LoU�����^snV������ѫ