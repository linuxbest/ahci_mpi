XlxV64EB    28bc     c00�ٖ��p�����߳ \��(~�b��C/3�Y���M�2	HV�� p�B�_���)��BCO@ݕ��;�I?ޠx�|w���w��9E��MtR�Xn���!�=���3$?̖��D���etZ�1�n��羚7���]g��X?4�Z|	4^����H�@���F������E�DM�6ԡB<pBxg1�Ɲ��Al��c�%eh�?5��@.S��קk�]��cۺ ���9�%��lR5��lr�0�g	6���@�_[���H���&��,��P�ף��@y�Ӎۍ�n��v<я����$N$��1��ݦ�I�X܃;PkG�lnΚ���P ���4�����)J jM���x=
s�g�����㲣��/��x�7K�sÓR��ܪ��KC�/�B�~�.G����q���v���x!択�ǯm���7�38qEP���@��m�A����&O4�Thh�3�Yv�I���x[�Q�
4�(�Fvݙ�Ǝs�Ӝ��ygU��d��똇"f��Fp����-nWS/хF�*kZҏ�^�~J'^�%�p`5��)!J��3�G�n���0�. s��_-��++D�X�Z�ʙ���N�"��E:�j��M<t	bA�i�_i�)Nr������	�2�D���#`��$e$�բ�Ǚ�0-[Ecv����]td�>y��1S<d�τ��~�����0	�����ýiFδk�bM���.}Ν�ƀ�-�!fL_�ۘ��l���$f>�Б�>l.\d����A( e3y��ڨ��l���|]�=��H����S������jo$�%z~:�:b�q�hy F\�)�H�v~�q*�d��C������6_$r�&�V��Y�VZ�W�C�f�Zia~.���Eh�
�ʉ�.Q���ܰ��Q��_.�YۡԜ�t�d�r�P-�҆��(5�z����{�<�ecAF�o|Zb�v [�RC�L��&�yK�i�]��3�G�v�"�z����Pw{����˰� w]������T��@��õq �_н7�a�@o��K��x����i��)��D���ꬁ�&诙ǁ�����{�bt�h4A�>
c�w�]ͲDG���X% �>��~���]��Ɛ<����S�s�T�}���Q$�Ǖ�3��i�<�r�+�2��%�Kk�e�H�I���F�yl�{�ӊ?n��[,DU�-{j�.ak����Ԕ���U#V]U�n� IbT�[����54�֔*|��*~�1�.��[L�۷�+�*�bS�ų9!�A�����Z�Y�L�u��9�{��w�Qb���(��I 2ٽSٟ��&�4�ӳD��ց������
�7�����8��CX��Z��)D ��}�D��3Zc.�S���<a��=sM�̬�,��$�2
۸�.�;:\�:��ݪQ��@�H��G�{")�3���.-������
�f�#�r���AP�֋
)��)��I>!�T�wLܾ��\v,F��D���`�����%�㞱L�_X��'p]��a��Lw�H���F���0��i�#��:΋�P��|�Zc��>b�i�`�>�^�@adǚ����1�t����3�俬�8�E�RtWHA s�>J^�벰mI�~	�
D{e�6�G?�t�W�|��#~�kߤb���,}���le�P�i_��\�����i#K=�nY��8�9���� ZH5k\X��tfv���hM*�x�m5�殢�Y	c6�̢62J���"���-���yS����}]9�֑͎���>j��m�H�wx���g#nܪ�w�x�SR`���dK_��e�&OOX��`�;Z�|�c%��a�*W������E�G\QE�na���j�Y�'m�X/>x�E�(?��̞�^�pE6����r��iK��Z��TЪ��
C���Ç����<�7�T�T�3©�]��h�B�k��;;֭ٟ�[�[Djx�ٽ8�TxS�p�\	+z6'�^�0xhzÐ�r�A�`�@0C_��u��y��
Wb�Z>���f�`�T:(��0��R� �qZ�>��:f�B_X���3/�z0�i����_�_�V�N4�^|��r��!)�#�%�B>mT��l��z��	�4��(�uv�����2����`Y�Ljk�{8B�h-�q7�kg\�B�:6,ɀ���WY��z���*Z��N�)|g
t��c�g�\�K4���ܣ�ۖg���bq�|�w����_���9ܝ>�&kR�&�D�_5 r�L71�/�����g���W�ຐH��ŗ�/P���8wvi�8��th��2bBK��c!�$���t�/ʝ�'#�-�X77�Μ�}^	�xb$;�K�3�3>t�9����.�֮\�$�a�/8�( n�e(Wd[9���h^�1�N�ε����T)�Z?آ%v �T���lb�i��L��N���i��� P"����2*ĖX8�w���q����6�_S���!���'Y��u�Q�Ƣ�^�A�iVe�Y�X��@�%�|u���&c��9@2P���ܮ01�Nf����0�^��:ԓ�E�Q;WB����!�)cTj�� �Z,�ՁQ5���mJ3
!��\��,�H  �����h�\�v��V\�G1�-��\��j˯�k�$�o�\~c;J!����]BYVk��"w�b&*���{n���R��!�j�V�i�v��Z��pp{�7J�Uӂ�짧�<�2u,�9�LD|o��n��;�.l'�k�͒�a���4@���s_��XD$���Ƅ?��B����/�D��+c�3s�҆���&���p�����������V��d�v�k�4f���QY#W~�E��ͅl�PLysЖ�2 W��p
�jq�4WP$�Z%��#��P�y��.&��It����!�ť0���=R�7�.S�����5�7)�6>䊇:	Gx��IQ��A��c�AX��|at���� ��%�=-���C�rpe��/�e�n�T�ݱ'o	��