XlxV64EB    73f2    1710-��������ؚ��2v�-�Ξ�����<�x	��q<���L,B.h�}w%/�J(��-�@�K>	�O��C�
+ �l~EY�"�2�Nő�栙xf�m��i�-��y�����.#�1��8�0��E����}57��N�ݯ㏚�U��f&X5v�8zh�gRj�u���ՏW�%��V(/B�O��巽����=��gQ`�����q�n����5m&ڪ,��O8������N��W��2�щ ;h�K�W���S3����^�4�a���G�>�e�#:�#M�K|�8~�p�6��f�P��L~ch[^����3Z� ~�%��>u:<!�e"-��GLb�nm����q�t~�(�|S��Tk�5i��'�n����*t��_JWo�k�C��ƾ�,�����M������KF&�ƃ<��b(�=!M��_ҽO廨QY�^��^|A��~}����^� q�	�����V8�<i���0��{0k+��T������C����.���鍋��̳���	��ԱLm]�Vz��TR=�9�T����K��S �I�S����]���iƺK}Z� �g�IU��r80cR�y�Sc˄أt��mW��{�?vR1����)x��.��r��˖PdҎ�Zu�a��Tܝ���Á����*��3�Z���r*50J�2�rR!I���S�������ւ�%��s8��Jq�i�JI�/4fǁ�ʿ���}����k(��vv�"�Dη�%Sr�4Q��ؐ �$��9���yε�%ˠ�wI��`/���]���E�7���.�3�60���yj�D~u:<ҙ��!;���h�E����G�N���D?	���O��8���;AJ���X>0M�87g;�
�F}v���w��
��A�Ϭ��)i*�9�J��_�l��y����
�GR��Mb����ZZ�S�w�$��l�Qv?��qj�OupY����[�eR�I�Uگ5�a���ێԞKԣ��s��Hj]��B]>�����8�"[m�̋�����!� q*�/8�Y���	�!��6龊r�Mٌ:$nƜ�w��,>���9[�o����z�F�~�81��I�4�Ni�9b�X��X��z@6��h��c���5%�W�-(C��yeܡhQ$�ď�ԕbZG��;Yt��%r�by=svd�jڅMIR�q�+4p$}j��QS�7~ئ$����j�?NYa|����|x5��U��+�_8�ic�',��Ys�g�W��|�_1�uv6�Uz�"if-��i�E�ٻlցV��J��J�-A�D�w�ȸĠ[up$�g@Y�w�4�D���м��Ǹ����
�d����N�?����\��WL��a�(B!���T qL���'���S�\����9,J��O^���G���A䕴C�Uw�췾e�M}�b)�︿T?f�R�]-���/3A�zH���'���c�>yJ=^���;N�4��86$�UV*-��FC�:���=.�[�/֜Em����%B�y�� ]�FFn�*}�(>�r-�)O ���Z��ލt=}��\j��v!�e}�#�C�>�P�7������}N�k*���2Ҙ�ưkA[tS��\��>4t<�K`�i�=��'Y��庑1/�z�E\��\���,vK��O1_%����m@!&���/�_�?K�(�	�Y�v���n�+�?�W��K<]�*���v�N�7U�$���o�G��fŃs�C�����OYi$4��P�z;�މ�����tz��!����
�7���-of�V���k�铇y��4�0 ��b����G ���S��$�SM�_�:���F!���\G$���11����L �ʩ]PvȏB7�(��(#����<�p�;���~RS;R�P���z�v~������=�]�ܧ�o�YTKq�0A�+<����#��c��6���<t��'��4��L4�+BE1}���e ��&kGϮM��� � �S0�T��$�D��0GH�4�H4��
�@���ͺW� &��7 �����齝��TDI���a��f��B����1�M����U�*�}�4���'�~w�I����D�0��V����*��O�& @ި���C&��)+��{p�X�C��܆ W��xŗ����6�y"Ƿqu�r���$�!x���"	Q�s]|a�]�N���-$�e��d��Ys�ϧp�+�8Hv	Qr������w�=�
����k��6�w�pk�z
.k6т�����ҫ?�>w';�8��p�Ǉ���@Nw3�oZ/�(�?��[�U�x3�GS��.a�	�,IX�
e�[T���U��~�bHE̾yۗ�h��e)��+�������7�B%KQQA�aC��Wɛ*���<;OOkU�A��4�.S�iM��}C�5�Y���z�9��ݍ���CDl�I��. K8�����H�ԁ �ξ�B% �� ��-RN���=��M�	��ࡓ�p*E�w)_vD�
���,�1q;jO��͌���/�z�$U�E0����n\�#r3�>"w����A����f��E�<��v[W�f���$��-���Z;J�A���^S�7��q�0�d� )�* ��x�>����L�r_��ӿ�݆C��y.:���O K_��/6�͊�2!2��(ƪu�ղ�YkA=�Ĳ����W�ﳉ��m�������3IL6��B��^ݼ)��|�ן�����G�J
<Ew�פ�r���	,K��v*��+ot�'G4&���`!����p��Õ��V�!:.JȆ�{Ɂa���g�Db��kJ�'O�	�,�1���?����}/���DF@3���{߷�����D�1ɛ;W�G��&�����0�����@ߢm����I��#���|�tQ�6�	3�Od��X���ӓ���-1��%�2\}��F�́������R��H)T(�Є!��G~�a�h�1������.DS�t��4@�10�92A<��Ʌ_�M�)�Z�{��������$ñF�����]�*�f���-�	���q���7|e��I_�Ur(��9U�X!�,�w�FD��愡'�0�s?Hh�{n�C��?��1��|o��f._Ե�j���뛡��̌��)�xƷ7߼�,���!�$�Q�
�^�G�]fv3�#�
Jm|�T��9�D0c��ڢ;��<C�&׌�FbqT#�*;z~���I�|�m)tI ��	\i�Μ ������,�٩�aE�P�+�,���q<�Ԥ�LEI���`�?�i��C��F�xt!�>3�W�[�>\^"�k�L�6�a�w	����p���Y�U4�tL������F�	&�F%�J͍�Ɩ�8�qRox����6���k����Χ�M	�>h�$9��?j�7>�r^�/��3T�z���->^xI��a5��F`�z��cJ����a0
��x.d����)�TD�>W�F���ca!V6@���[(Wqs�I �^ՠ;1T��� �n�S��������H������{�� ˁ���u7U�Xv���EE~�,[n^�� �O��fB=_�T���2I�;*��U!�>d�N�:�ln?��y�.?��	��6�S���g��n{0���l�7k�䢗VA��m:�ôhk�}��i��r*J篜P���5�iÛ�a��$?z8��AV#7}�`* 
�l�@E!&ݝ�[`�)4���szDɩ�(�NR>r,l�c/dv��(bG�����G����d㻽[uZ}}NE����m�ʓ 	�Y?�T�I�D��ʛ���4<���	��Pg��@`���x��d6��'s������V:44F��'�	8n���$�2F�DXIA�[�����6��X�W���Q��{X#���h����t�n.n�0Re���t��[���To�Cf�ʷ7f��ny5��U,��$첹�\'�.�������0_#�	���```���{6����ĐWm�4V�ֳ�9[�~����^nU���?
M0|��z��`������&=��hL��KK{�a��;=g(�j�_]��@V9sg�����5wԏ�-�s���qǐ�N��J��lq�b}��5��D��Q=�g�98h�O���]=�%z`6�3*��Y�TnHѽ�-�T��	/Z��t]�rʫ�,)x�)B\���3��b����汋�ݮ��乣�2r���n.��6W�H��,�Qxvr��4�ki�Y-_�.k;� �]G�w�jH�^`�i�/ sm�$� �2L�-�3��JcaN��0���-/}F�׋)��!�CDK��)f#��]�'X��_5�<�XԢg�M�L��"�<��J����_}$.��Qd薥�FϡK
�T�֞t��ɕ�{��R�J����E��%`��v:��*������)�_[8�`���O��Y�9 ��	�61Yv��4��l��������N�9J�ͣ&=�JYlp�w�T3Q���TIuX�Cpࡤ
�f3�"![%�:g�c���ޥ������B9v��MU�<�0/Aǥ�~$Ġ��l 6k��zw�j���:��k���*��5g�"S�εx8<�v(l�(.1T&���x
R�f/>�v���`;�,��R���q�2��|>��{��,����IBs�)ùpL�^�:V��M}��W��_�j�i��TVܽ�V�~j����6�Շ��c5@h��T��Te��L�������g:G��m�����	�:��"^����8P4���wG,�^���@����A�J}�G&,c���.D3�|恜���&�|=?�/�a0�Q�,��{�|gm���A�P��sp�<�o� ,��p'����qr�����73��{��sw�\!`���#��ᄋP����9�n��*�"�Z�0Xw�p',���|􀮮>�>@�`DޚN��iJDv�p��[��U���n�B�A�LXSe�B��x���[#Q�ȴ�g��ӎpD�E��]7�7̽�}B*�t�p�.�� �[�´o+��ăAS~?~4;c���31]��:��޽�I4ڳ[lH��B��n���i���?�g��}�+r���X&���K�K�̘�(�Q�iE���x�ղ�Iv��sm&�`���}a��TH��b�HI;���� 
���Ԗ��2'�E f�{$����ȕ�TeM�s*B�ތ��8����P�� �b���k����\,­��`�;T䄫�͌.fwF���/n�f�^�h�b������q�5a����u�2)~�T.40vWus�th�2r�~�d��G�L��!H�'��V�� ÎBc"�֔F���I�l���2u� ���4$/9�N��j-n��+�������H�O��A�Utqe;�.GWx�%!��P���_�[]Y_l�(}���	���|��'��*tߗ���o�N0�����g X��'!WLd��ocɣ!�|�xO��֓�� ������1��z�v�1�i쟬iW�(z�_�em օ�XwNݵ�r�An@+X1���q���KX��.��� 	�o����i`@bEx6�.���ђ��֎<�~Q�⩘��]I�a�%��<��%)~Cd�8KSsi􇳼��W�"ɍ�^��1.�fCEZ����"4 �2�K��P��"��#HYbQ��t������rC��
�%��+l�p/���\ �mL�'�c#�J�8lL��d:�Q�#���`n�������
��Z ��P%����j�`Ydb0>�$��C��;HE�S�[̪d�ޭ�",�0����