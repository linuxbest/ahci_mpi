XlxV64EB    fa00    30a0r�P����Cx<��pS�O?RruN}u���"m�Þ9؎/�~��}�Q�W���F��fyD��
P"0.N�s�喉��A�m��3�M�U�_�:'e��2�8p���G�L;n�7�c����#�x��T���^8��}��}���W��Oi�I��3X�j`����*��q��'[������N���0�tt@�ކb�E�K�<���C�eC���ND@���@D�n�#�t)6�0)���quh��6q�W��_�#���Ah��L�4����q�iQ�E�m|_y
�^�W��+ [!\Gv�v�;u�
��HgR{�2CАA;kn|<$�%Xl�X�C!J�K�"��(�ޙ�Z��Z�HJ�m}��·���bP�=�>��kb����+�(���H5���C��1p�ƌ�3�ua�F�ˬb�0��,��g�h���I�s��9��஘;Þ��du�'��\�@Z�z+C����S�nH�?��bƲکS}�r��W����.��c��5%?�p�
���̫҅`?�qd�[��C��F��S�Gچ*�8���5�9 �-���W�.oea2t��>�R� �0���5���~�<(�8֤ �u_�U𭶘�i�,���E��h��!ϙ��B�� Ь=Fb�$�U�S2>[�bg�7e�S�?�mQ�U��5I�y�Y#n
��䃥"� ��%��z�j�&��S"vy��C`ɉBr!��	�c��yضKXRQ�]W��m�`Sn��Uw��ǥ���D|\G��|0❹��u/���Dt�yL����,�V]�|ølq�$��iOb�!ھ��CRb���U�Kv���GL��O5���Es��Lќ/#,V�a8>�D��)�N$��/5h9��Ԡw�oИ����Q�<g;Y�,��0~��[[�����_�,���v���J��z�\��񵄪��Ւ�J[�r�&�٠����*ep��AW ��%I�i��h�l���S�2�\�,
p�$� /����V���8[���zL#WC���r�����,�H�1{�k1e�'���<W|��m�*�9`O�n&s�˞x%@j��kk2����h���Ȍ�c������	^4{�[����B�E�h$������ͯ>V��֑-AB��6x��z&K��7�+�	��K�ԛ40M��*�� R�b�ب%�O
���H�M�W	8|��%�͡�0�˿Q>xj�jq��~ L���IU�Y66�����xsO�{��E��S��?����� �}W��C�?�����'���(�ϱ��s����\���j�t�_^K	���yOg�z/��Ѝ.-7҄���o%�Ǻqn<Z=�U�g�,֜�)c��7TNlDO���ev�qL��&gh�MP��@m����T��%M��a�0��㼅9N `yd�}C��B��n��vy Tgé��]C��OGdx[��h�%���2Uʠ��X��|��m~�������ֿW�oX�Z���Y����Q#~�D�{;'��g�Q�����<�r�ޚ�e���������pV%�%��B��>�?��|*�e���C���Ub`��,ظ [�Y��d�.A%���#
��Kp��< �ͷ7_����	��a��:�A�u�DsD~w�#+p���-��K'N �T��.9ĻQ����NMk�s�i�)X��6K�8g���v��t����8cLPFg)�N�t}9��.:����
T_��FVV�x�� ����a��9�2)G���Oɶ� �0�%Ǵ$��CA��������2��ރ�3��w	�S����L�]�yR�q�WO<��[Xj<EU���OU����?���6K�,�\B�A����nF�I~"�袅y��c�%W;b,Yc+�l�H�4ԉϩ��K��5l�Fj�wA��
C�t/�ْJ�"\<'���� �R����7�Z��!�U�GBv�I[�������.����	ʠr��⃣�b�|_�*��D"�b{�e�ΙyJ��g��-�)��.����5ڑ�-yTV�3\���;<��n�s�.��#�l?�غ6�k���#�e<�]g%��w��I�E�}^bF���;��}��XQ���(�e.)��ؐ��@�|>�9>���/|;���T �$Ga�T���,��74:�;5_udC��5AwCJ�3��FG�O7����6�k��+7d��@����/q@�;�蒐�s�������GFr	���@J�y[i8�[�E�G�Y�X�<x^A`Y��4i�HX h���L���� ��->�� �G��+J��4���f�eڣ��]K�ܓߗ��~����.B��Ja����V�s�x����nk��p��T"[d��|O���j,P���hQ��(d�u�g_�3�]�I)mK��ױ���&�5��-�]t�ũם����>�>�����@�Œ(��\��8讟��Y��a����1���.z)	DM�y,·%���?�t� ���}����7�sl��E�����&�۩ӱk��2��N�d��xS��7�o���i�,�oL��#��z�
Z����!�[�"� ���~��(�D��!Q,d��$ �)��"ny�{�}:s�x�wz�o�b ��?6o�v�	��@v�]��%��>W5�Q���j1�39h����r8�]�|����UȎj��IO��Uv�?�TK���p��;z 6�q�E��?��o)��� ˪��xEk_@���X�2ݳa�ү%$��Xn|QIH8��q���D���>�Q�?��oEKg��w\q4��2#ɡ���P�I�+	�QKOq��D���8�E�b����˭���|���Ox��b���
%��*�dFu��[�u����iQ��ٜjuH�Hy�N ��s�@xɍ�[�����ީ�s1�6�kZ*صF QȗyI�_Δ��S�ɖt�|�}�,Qb�Zcj�*7N5:��{��q�'�ݧ�E�1#���|�l��Mm���*�'�$��S�Z�Nz���^���`��1��.W6��U��5��Z@f�ˡ�$���Y��9xy�d�+�y���U, ��̴�-!ό�������h�w�~�E�v�^������o��j#���(7ߋ��E��H:L�G�$���:��(%�����vC�Ǚ�r4z��]"�{���G�,{�D1-��Ё�>6��D���gE�y.�W�M692�3f���|(��Tz]c��a^�����z<����SrP,%�����5+�&�z��i�\ � �Ȯ�T��/q(c�쇉@��BP ���߷��^%�/[���-�@l���2�_tKB|k�:V��b�	�:�5w��Y���v�$ۖܢT7H�C�+5�9\i���7��3��NRc�9X|�BȜ�(y ��.��/���C�����㢐�l�)�hQ�����_��ʭ�ډj�k�� iL���R�ؐ�gxu�Z�v�B���q��h��_B�g�+�߳����mY�(��j��Kn�Ղ�kœ��Z/�Z�Tnc/��"��{��G�5��,&ޓm-���v��L�/��A���)�.�K�Lg�x	$�PJFY�Nj��V��-p�嵥Ʌx"�`!&��� ӎ��פ3�����W%��K���T�OX�tOn)���Ou�p�Y��(謇%�:���.�Ͻ7��#O�ﰐ<!UeGE�������j�f��k�)s.u�~�����F�u0<�������$0�_�y��6m�����Sv��JŪ��ʳ�����.�b�"x���[s�GB��x%~��s���������"*��p�8���>qOl*ǭ��f�c=�[Ԩ�����p�6�ZH����y­s��ݔ���J��YY���>�e��|ӥϖ�`s�u��N׼5v�	<{U����A{B0M�t1W�ZD�I�}���P=Ju?'�e@�N�#9�xAS��Rg���Sf��j3�#�T�Z��������7;������F�*��*���{$��0P���L�G���.	R�l��C�T�eh��:<(��/:CD��؊�f�j8�U��lRJ%��虀�R��2U��Tt׎g���$s���e�&8� �W�鶆D���F���~���n��O�>2 �$,�v��7�h�F�*�Y���?�	G~i��x�BE�48-������9�(����u#�M��_)1ʹL�O�X[���\5碰jت���^!*�1�t�����A��f�C�k��Aw�;䠁�[��8x&[>��w4���^1���3���ޱw�<���X�r�hH8~t����qȼ����;��e��~Sm�!;}��a:e�z�/�jU5��i�J�������o�EBC�B3%E���$ ���yp�	y4�ZP�-��r����1i�"!�#�!9�HaŴ6g)L(�(�7@'Jѯ�_�~�R���g��
$3�(��ӐS���9#��F+tQ���\����' �}�|���ݴ#>��q,3�<7��5�˂d��_j��QJ_�xГ��@Yі��Z^���Yb�����tM.E�Q�ԂX��6��^��n'�5H|����ם�d��c�U�k�e�^���ď�bC9�OQek�`6vڏ�Ad��9�p����զVG��҂������1�xz�K���%�V]��`ٟ3��(cx�0����R<��U���TzH)&�@ 
�ʱlN:�؛k�ݩ����@��\��T?:��>.g�(�o{�s��%ΠQ@�E�v=�������"c�A�`7�y}F����x��z�d���h��T�I�F	~n�C�	���
�ʄ���C1�Bc����~�m���p��K�k ��(��
��P����p�:�ȸ�g�`_ �z��8v��2� �.��k��+��A�ޜ�ɕ
�X��4�M�%��'V��NS�W[F<��
G�?2J�
uRS���z$�����ʆ��V%�d�����F}=�{��ZI�=eO�����
���o��W���
u$`�$ $y�&��?��Ғl�c�L�t��?N���m_L߄�1�P�����#h[dI���+�?�A=|N�#����3��c��q�xC��Q�j,N-��lMb��Bۈ/�����B�?�=�$ۜ�1�f�սQ�l3���33{s'l\̵�k�Îm�@T��/<��*�����5X'Ԡ�$�C��ȯ�������$tb�m�U;�#G�6�@*OE�$�z��u����Qq�6�y�D�9�-��׈��0Ȅ�iL;N�;"� Ԙ�c~t��M7�p��� '�v$2�D�rE������+ m�r,��}"�@�{�,oy�����������·.K�	0���d��q��;s?��Q.RQ�����
�u���D�����<�PX�}�I��!mG!���]`*Ѳ�����/o]�>ѱ��AJ ���zľY�ƛ����W�A�}�k�E�QZ�2�eU�W/�}��,m,ᝉ�*a��=�¶i���'d=�H����F牫������� ΀�ѿ,K�S"���ԑl�nP��Ϯ�Z3|�B7o����e��{�Q��e��eѦ��Õ3~nT�� ��B[˥UN�V�f�&On��	�N���钄�4���hxJJm��HO�:�]��AB��׌ Ǯ�2u�S���3Ꙓ)5sq������Yx��E�ԨLq�&&; {���G�X�*�����) ScV �,������ E"���c���0F�t��b��N�b���H�?j�D��r.�j����-ZB���о�;g )A�N�GD���#�w0M�|`�3��g��?ު'�����T���tN@�yg��F��ߓ��&g��)�b���=�.:ӎve�3F��9�Bm��Ue�t���:�6VnT�cނ�%�/ u�(��h��|�*�˵�E��H����V�<Y�Sq���	0#�Z�B0Y�$�'W�y���'<��6�����w�Z�iT�s��ZS�0?�ݲ�8K✹}v�"^ A��2޶�Z�F���~ps�8U^�$)�H~�af��n�aZ��8�
�<��{�����I��\=�fM)M~���9�)�����	��41��*A)�bԼ�� �<!�w'���*�z#vɎ RlnZ�u�;"9SP~�<�q�l���ւ����d�=��I�#����y�XX~�\������m������ �\��C�� ڶ*{�y�ΣN3lqXUG뺠�i�8ׂ���Z�w��}5���"��+^�Y�u�0�ӆC�Rvt�����)���q����L�:8��~�d��$�x^R"l���S�\�L]��1�E]ue�؝%֭�[,�� Q�����5[#2�毾�؉:/��-�sb*'I�)��l㐭�g?�bo1��� ��8��5	�urW�8�k�A�����z�JF���<V,�����L�}u�Ԫ�l��꡴��:ؖ#'(P�w�<����I�G��Y��Ě��e��hS K�����l�p����؛w�����˩KT�75w���\Wϡ�^I0�Q�ՓȲ��5'�8��6I�&_���򵽄c�Ŵ?ɴ��8���'ڃA�%��O���Z�I]@����j��q���N�=\�S#�q9x<����~I�Ǒ�j����(�t@�z��B V�Uk�蜒3)�_9�~rD���x��H����?ǞyJ'�����g��͖���j+�5ک����p��z�8���<�D�(��}
�*��}x��U�!�3����Gv�K�\�~V�^ҳ�.�ﲲY�V>i��+���D?���6��f�l�d�Kw���J�A8$�_;b�v�jeHIL"����$܉ɪd��J�÷�!�e����?���<���P2���Qt�r��`����ƅ$.*@��qT�,Y�#B�����T�� ��xv*���x��b�r��z��Ud��e�����.�Cx/�&u�a���u(3�~�_�?��_^���>���ň��i��{~��暎����q����H/�荲n�V�H4�Ԅs;��2P����^G6:6+���P���!K�7��	*�c%˝ѿ�*�>�c�xvk��C��l�8ӏ�r�u�Ǫ�qO�~D
g)P�[�~��g}nV�u�����H�b�5����@й�컒�9��k���L��`j|�č���U��l7�q*��y3�ޞL�be�(�(���������#�yf�5�����S��`2���s�8��G"Rl���d��ܵ�S-� �:�����}�|\��2d���ۗk)� d��ȘҦC���{����r��0�K�g�rHl�O�8��A���o�Ϙ���7w���4�	���r��RLl�zc�p�6k��ga �:e^����BD�̮��$C[��̒�yX��.x��< ���-�ݖ)���I:�Q��C�{-����IZ�2�j��W7����D`�*�%�� JXWa�� e�u��u��/)���b�|*�g^o��F+m�����=z�m^*�����xl֝�(Y0EU��b��hQ���Zt���n�%���"a��J�ud�c�����{�l�⿖��Nh�r���L3� Æ�upl�����ـ�p���+��U�NHU��V?�m)S�
n����1�5�i��M~{3si$c��{�z�l�FV�32��j0�3c�Z�8�.w���}�$�Y��;��{��	Z�",���J�Ĺ\ф�	;`�]H�\��5T�kT��'�w�E��Xp����C��?���m<ă��jј!�d�k�@>]x�	�����v ǧW�y�F���}I:�a�P�N���O���C����F���`ߏ���FP=حOv��oX=���/|�����'��c����t��LZn$�n���ЄC(a#VбyA�:K>KM�w�q�κ�&B�qX�y��MY�	���,�}�t醀�4���J�'�����0	����F�
q�%dSw9���R-�����#h��y-��:����.Vg�=Y��S7�K�q�"]!���y h���hR��g���`�V�!϶¦�ڎ��	ڣ��Z~`z! !�+"���~-��7s�ӝ�,���8�+e�X�A�X�n�W;N�'��;�I�%�?�����&^�ޫBwQ�Y^�����һe���~�5v��O�$��Ҹ�����һm{3�5����K��;/]1��X���p3����bϸ�/k�]����I�>�,+ ���E�y��D�wj�C�÷����\?7̶�*/"#[��,��:,lI@�pC�{bPK��� ��z�s���{� /*����f�S7ʄ�揫�0G�P/��a��f��񕂯I;n�;O�Ϙ�W�XQTy����H��� E���[�I�DO'�_-�I�!q�2��/���Lc��],��h�:wV���s~��>0����Z_|�<z|����+�lP�pI��%k޺.����r����o�eMFdQ�M��.�����	al6?
оΆ�����y�>�����͇6(��_>���a ]�_!uR� j"�{ ̙}�^����Hq/��e��#�L#��8���l�J`eb�� �gW8u-C�a�"���#æw{ �����)]Xx_�&u� � ވ��sLͨy�n�ߪ�:_Ǡܖ�j&M��|�_7�Udܩ�C���^-MS.�5�D���>�PA��^?1\!�-��{/�]�������cZ_y5�O���>xhsi�+q�w�Q\��Ic�#�.�����qyE|��]��}2U$�
V�h7'���n�BۆRG��SQ�F~�h�b��[�-����$Ԫ#��S���sk���^M�'��E7׃{���n�\&z�� �`�7mRS�M�@YG�e��5�:��Vʻ��p`���-o2��U�{�VMo��ۉKj��0l���F�7�`_�P�<�rǉ���7{�� ���*hA�pt�1%�أp�z�G�6
�$%�Yܿ^��qxLƠ��H�s~��V�)i\[��H�>Vz�M���F����\��n̺�R�z�}�%���%��t�'AO�..閯����$��iWw�h�)��C�#�BM����mW�������]�?����۾Nc�cxO�BS��^2��c̭x���o�#�0�����'��K�ii���Ȼ���ȀƟ��]��	��3���]�H;c�a�0.�y[]Q��<<jz��OH��|NA�Y����鵽�{9��l �{����վ�L��j*cg��Zqj�>��$g�n��Ε�ǓB�����޼fҤ2����႘��nk[�%���?��e'�4ɘP1p�}���LR7��L,rwj*��&�� ���rH�	)�Wأ��`a�J��"WF��TG��o�p�@���>^
j^�͆�Nc�>o܁M޹�F~��
�@ e|W�*��ׯ�%�uŞ���Y[��>UY����5�<�M�G���F�gc#��v\�ܻM�b������`̚1�WO���8У*5�X�sdS��wRAcs�8I�|���:o�դ+k�(�z�}wR�'s��~:��*X�,�h޷�3A��-�w��8�ؑ0���m�T$��͔�nw"]�<.��%���l�?�7���'�y� ��{"I�!���g�+���u�PKjE�$�ߐ���):�GI�R�V������_��n��M��7��dU܎s~�A ꨉV�g$�9J�w[�Ĉ�+@��g�ζU����Ʊ���aۢ�'`c��1.z�QE��S_"�,	ACn��~�ԣ�8T��')-��]���NŤ�t�l:�
�,�s� [���9is۶��0���u6q�#:�kO��[��D��g�/I'��@��{�;ł�h�ȍ���yo܏K�K�i�7c�"DyQ�ɋ���1���L��l;�_�[gB	��D/��8V�t[�K��l���68����$�W���.��&���?�ѝ�{d�D�ěy_y�V��c��)�� n�9�\�������z:yW��2\)�^	S��5����>�g�)p����cQlK��=��4���|<F��tK�BtNs�����'3P��-)`1�Y5 Ό�� ���\u1O��S��~,�f����Ƿ���(~�3im��B͟S��?��S)N%B}0R��9�ͣ�=D0:�0�17.W�µ%�vw�K���L��崢��(r�ا��؀.;� )n���VDODO^�9�W����J�Y���#��y(�	y�1֌4��.���!QH��RL�b�f�(����e�2�̊�X�̐nK���Q$���5��g�e�}�*^l��4��svI!F������;'�C���+��6���<�����;A�<k%�aO�K!N��z}X�GlC����tV���^��/Y3\Ţ��j��߇r?�kW��!if�N��ׯS~��k�33�ɂo앩T
[ʹA�o�Vgd6x�81W�u�܇�6�M_`'\x�(% ^��b{d�b��(-H��=�7�rM������~<���^0$�oFT>�	^ ��k�%I���D�cO ErX�I�8Ş��Ũ�١����J���>m�4<K������������R�	�t��?i+S�j7�V�w�^XvM�
�������}�c�}=�B�Z��sV�rE(��R
�I����,UD�~�jwp^���"$M�b�mv�-���>�}�H:s� k35fa1Վ,��No��5�)$:�,�Z�7	,������*�C���+\]Vr0m3Ti��A�W��V�P��O�R4鲸PF��]k��0
��8B`:0�5)�I�ܿ��C�^^�-S��SZ�4J�L�lg�5�r�;�an�����_WpCnu6>^OG�^���/�qH��şP=��>� ��d�6���n5@Xb�`"��1$����=��%��~ ιA� �I�}@ȲCzX��6�i���,<2ǟ?��m-�	����w�h�o���߸[�ek:�>ϲ>C��^���Ŵl�9�r=���nO�����30:7�0��0/Ϫ��"��&c��;����_�/�Z�SRKi�����dj�j��{h�A�	�����,ͭ� $�.ϑ\����c5�ư��w@�Ʌ�į�╮X���Ӥ�|���Q�֍�np�eTc>�y�E�fyD˯N�����M���@k�Ca�z�� Dkj<5o�y~n)N鑯����R[�Pg��g�XV!�"6�鹏�^J7nw4�/��r��O��dR:2�!�N-j�[�)F�by*��X����{�D;ъ��_h���D�
lĲ�m&� �$LZxl��P���.~���'é����Xo_C��|CR�'rbᜐ��1�����V��X���/=���ڇu%����&����x%��L�-I�đ��t�|�����Z�E�������3G"B�ԢO�J�9�J2���]�D���ܦt���/����%�����Y�a�<C�,,��8�4�� �
/>�J���3m��S�|�(���Z1�=�z��'���uM���M6�quY]N�M�|��]_\���D}���]�5���S��"�[�ae�F4�k��A����-��r�����Ȍ��f�G4�M%��K*Y������!����N�ճ�ϒ�w��!q�,!��FE6�����/H�jť��.��-J���U}��\x!�?�\�0�M��`'�����x�T�742�*fI�j��o�=z���cS	���X�wl/2KW���Dx��n4�6`0o�}��Ovԉ:�7��?�1���4�7���UL�͕VL�v�t�%<�fcIq�h���j�����q�1�Ku���SEAN3���`�a������	љ;��\uec|��H�:z��L0�����iY�Wܱ��ܮ%wU�U��2+�W�X��ϑ����N�2|��Zx���\{��w��.A��#?렏~ާ�(lo]�g��dWu͙@�`D/�usp�&�EvU�xxa�^wX$�2�pX�
-bJ�E"1�ˬ�a� �x�S��,�&�����b2�}����v�^�u�N�k6�e��c�퐙��ݯ�?u��4�m���B[�n¼�����XRiئ,����c�F�p�$��\Տ4Q;�6m���	9�:���@i2I�8W#n w���(	p8��w��)��q_�lU,��+�1w�����p	��5�y�#�����}�V�BZd�4���tu�ZĀ42IȾ� 'l�.�2�a;�[���&1�H�'9�������te�=X���({�v,��sh�XlxV64EB    fa00    2ba0ݷ'4TrE�-�L��K�b�e�Q��J�]��/)�ڜ����Q�%�:'��/��_ϑ�ԗ���?3!���M�w*��@��^%��N�xC�ܫ���l��wgL`5���$��d������8-d#�gT 8�r��$�����l�t p�>O����	d ��*�C�C���̶�U�`X�۵}f�I��9���R
�1�w����7ϴ��@}�mP/�b����Y����an�I	�~�a#i,��)��N���ߕ :_���W���o�?C����|)*AǑ�p��S�W&�>����E��;Bw� ��ϐYdn��ht�tbhI���2c��:����F墶x�Q'�7��)F|��(>9�;��_�0�ș�~�`��g�����6gj��[�̩!(�?;>���n0_8�f�ClA��#���F�	 ~VO�O���t"@��K��q�1jg�u����z5X��l��$��ٶ���fGx��-��b�Ο�ߏ-'��_�ځ���z�/k�p��m���j��HB��"��/��I��A���T��*`��o0�O�l(zJJ��A^5���'�:j�ѳ%���>h�������8�Yy��3,Z�m
�R-�%���oQe��]U�u'�i���+㴊�Q�H��?��2A�)��=;U#�Z*����
Kkؓ��*����^)���	�\¶i�>L�
�|��j�]L�d����}�5{��z#�4iS���/��+G��!z�R��ӡ��h[Iso&ޒ5�r�������"��A����
�(��(�n��PiON�ң�����6���ȇp�!���Q��ѣI!�5}m����l������{.��1?�Y}I�|h
]�i*�b�1�p=�������MC,�!��6��O+ڙ�t^;.�(c>w1��s)����xY���[�,l�fxH�r�r��-�tsi��	^ӹ~sg�c�ʏ�{3C��)0�^A�m����h�8C���J|r����?�1�8S����ɨ�{���B=H�X(X�����5�7ukxFU�bUZ�F̪�m�G��g��%�5��;��һ�~�+���l���|�2�`\|s��M��R�`ڮj��1�����E=eR,�%�/�P3ٍ���ʿ����n����Cl(�=��ȵ�A�]RD��ìjHP�]��%�'�.l��r����|��0�� T��UCl����F�Cb5{P�u��ݼ0���/ᬓ|'t�c�{���)�tP#/�X8ղ�IR��)������1-�����YM�FcM|��|F��Z5�c5%�1�J�ǗkY9h ����wp���#�)?��i�JR�l�Q,m/�kb�����Kխ	lg���gJ�#�b��Fs������{�m0����< �qX�Z &�S�X2��Q�@4��I���ۓ���<��sK2?���|�z�x$V���	`�����}��.L���D�=�[���C��畞]�~L�W��6c �����M'X8��Hi���\��VC@Z��ʝ�z��/C�ă���`4l3���E��#����2��,>�n��r{C�kzc��Ka����p�ǣD�.���ǔ"y�	�s�j��pT~�R�K��ğ(}5S��P�t��X_x�����р�m��HրV���2t�)�vYr^��p�XzM2���&5J�/z�#I17%|�f��Kiq`I���l�����^�u2Ft��M��Q�K�J>�о��h�
$oV����M���K|�3N;��(�}|�>�s���87�p��F��y��@���;��Q�[k����bJt���8>�k�R�Xwuv{]�"'�C�`ƅ�����T�����dEY�{3Z�G�b�Ϛ��F<�$%�C��,/?��R7��2#���F�lʚۻ0��"U��b�.b{�q��D�)(?p�1�H���UXn�b����91�)$�ϰ!�Ềv��s���~�e�K�K��K�F��`�t�&=����D9�6mg$�X8n�f8������!l���=��y<�aˏ@��Q8rA`9 a|���� ݵ6@m�p��a�FI�����y�H���\��]Aǉ���2��������W(k��c�To��a�u*����4�7[�7?� �(~�C�f��qpg;ք��f�b���j�X�H�g�y��g4��O/� ��ѓ��<~�dt�Z�Cև�{���.h�l����td�2���N�?!ɇI��f��������_F��$��a�F7"^H����P"[,M���c�0z>��3hJ�j�,��1v��_��*`�3u��x,i�?�߃1��s���4�U0$�UOĕ��	�Y��p^��i	̓7�6FBU.�>F�:�����N��ll:k?��d���v�ΔgYZ�.�KT�π�}�m�#���`
��q��k(v�2L`Y5�h[�Y�H������|P6)5�h���+6L����F�]�Cz{���ݸ�H����v�:��]wDς����z  H��s^1�wP�B���J,+��Z���ͼ�Ґ0���f���\u�}D%��l'F�hB6��Z���?T�
�S�
q�$��Yu�B,ecU��͛��`�%_��:\w�\}儇����uA�o�
����m��Qd�1y^���4��l
Hr��U�n�f�6&���I�D��v�w˗g���,�n�}����6#�G��'R�n�i�O2=����#
���;Ct�`�P� "&끆d�:����^��UxKs_F�P��3�Fv�]�
`�V�6�Ǒ�w�o'��C����.!R8����(��~��L]�/����i!�|I�*٨5Xr�0Y�J�4V6|����Q��ܨ�&�2���D���0%bi}�(s���YASX�6�ZLbY';/k�
����(�ڴ1�)m�h�"w}t�~�����#�#�"�׀Q1���͠��vp��ə8�֘B��72�:��B����B�r&u���my^`��!��1A}��Mb�X�[�� ��<|X��?���`�b�SQwsx������k.�EN��#~)q߉W.yn#uEA�:cI�(�_7lx���Зal%HF=�gB��A�3E�3������\gB�3bҦ^�ɪ{����v� 1�	���-'��c`�e Ѯ-u����a���̑.��W0+d1#��t9l��Im��T��bqN���-�~.P�h� �qR ol���͖�v���(0&Z h<�:/)��S��b�i���6᭾B<��ځ���U���|��#ȁ�d'<��,U���ؘ>E���Q�n]L&_������}���:)M=B��iW�@���� *xy� ]�|b���FA��g��	�I+�Q�-ڋ;���}�9��_�/�ڲ�"0��V�b���SC�~�j=�+� bx�jD䫙=�Þ���6�����@S,%;y�K+E;��滛������;���; ��
�JE�}�������D
2 �}*{V��\T|��{;�0/�U'�T�c,ɃM;M��o�D����!p<�
i����	����O��!'�o�m2ll��K���t��{�W�}��WlMC�,;�Rh�dH�w�C.����´���0���x���]�<C(}'�5*u/R�?�Be�ˡ��*����1����9+���	t�_��n�Xb�%9���Qe����a�OU��������\�N�[y۴�cu7���I���*�X׏݆���JR1���\?�GV��8N�U?iS*�&�$��e(W���hI�ƕdgPܷ-��.�eK���J�{�]�p��Se���k��fgw:��%
U�ر�D�+�/+��b��Q+S�����E�cڠgI�:1�Ӿ���� ��e ��L�^T�]ME�2�����t����F��:uÙDC���i�����2j���>�lS�r��0�lܡ��"k:L �&��mǏ�EFm�D9���=	g,Cc��rQa0W>���8j̱�����:��k�#�B�3�j�O ������r�
&��]�sx�-��%���r�n_+ƸP)g�f/���$&<��hƈa;o28�H}4���/\&k�y']��\��S���c�ۀ���r���O9	:���uZ/D%&v�3G#��$�W\%��q&�5�5�>5���̶R������2����?b9<e�%<1�]Գ�҈�֧�a<����H+.Ϫ�Xe��-F}T�	^��g F"�Uho��\ �1��m'YY%��kz�YK*)��l�l��+8����3Q^Β�'Nr|�+v�lt'���:��X��b4���@D�����ϐ�0i�u�1�Cd���߉����0e�
U�T���p�#��~M�� 21D}���9��w�P�ݔT^_�o�+���NZuz�}�V���֫�";ʛ� �r)N��+�'�i�9ߎW{ }Մ9��sl楧k��B�6+~NU����7�m']��7����B-���>�%���i�4i) [}�KU��Z��Z����ɐ�iQZ\� ���>�r󃊀C`�BENoCe8�Y��G/�}�A{,�	�	�^`�?��ozC��o����/9��
Hn50����6���B�b�|"�C����C\�ch�
'�n�y)���إ�w$�׋�w�lmhS�ƃ�q'�8y�f�M�Y-�@�sB�q����|O^qiQH���~�I��q��Nxe�-:��J}�`
P('��j)�%�JΊk���b���i����7������A鴯��������y���O��>>��l��j|���j;���.#l��9T���Y�B�q�����U�+:�S�,���쭱m��q���d;m�]�t!��Z�U������ή��YCJ����q�����'cK	�oL��]}�R��N�E�=��I��3�̩�j���/Zp�y�y���������a/��xˤ�vs��s$X/����F�y��^�g��ȑ�Z>����|��	%4�x]X�_��ؔ�arMiWχ@�^�w�|����5����1[Y�����K�7������ߠ�y��S�����Gd���:q���A:Z��[�,n��s�W=�z��T�veb�6���`7�Y}b��&
T�dv�8�v��i�E�$7���ׂ&�I&�b��&c���"B÷���5m����hY-�9#��YDI4��.b޳&>]�t��F�C�*C���q�p�xE�y���^�����g����\ �����Z����S���k�R_Cs�uHKj�� d]>�
$��!�1N���7��F�?���� ���ΐHٵm ��-��r����&��\��0UX++��,�#�Q`$�)�+O�u���0�����B�^��/XG���！ī�4`�ccqL�D�%��E� �<��YqGU.�'9ʡ�բ����7����c;�[9W�S�L{΋�VJ���`�ze������B�*��G����6�Ϭ(����,�ݰ�(wX

�L�`"?��� e/�U�Z��{��-y���&�0j�6wu=HRG�Mǃ�y���1�ݨ���c���]��߂��2��T�����`ɾ���1
�#$$\���-)A�|�7*i�J^�/Z��Q�-f��MK?���(�@u�J>�=0�ǑȨA_��p�ą�7kHf)D��E
Ғ�ӟ1��S)�<d�o6YO�f��,�Ũ��޺��=���%�y�Z�������9�*Kt(��c�1?�u�'+qPT믟���v�٦�,��#^���`�Ŵ��&�ێ{H��{�����]8z��*$�"o�P�p����g�2,�8��GN�rn�� #l���Z�E����x��\.Q��iE�鰭��&9��	�[ᗪa�uLe��p�W얭;�!Q})���|�N5ޙ\�c<�ş��͡�?e��wl�2��L�7J~D�A�і\j@>;d�F�᦬�&9)���0�n���]	�H��9�*�kHv�K��
w!`]'ݦ���}?x������e;'�<ݗ� 
�a���'�E���)��]&sBq,D��?����;���	��b�}1=VQ��o�c�B:s%�q�N��A`��N1�!X�7��e1@���	ƈ�bT1/+��mS>'��^D^9r��A�MG)%[l�j?0_�eəG��ز�6Q��J�E�'�4��۷7��)�7��+s�45�9��]���t� 1#���W�<�0��k�Y�;��0,���Б�W{;���\,�"%(�_�̎?ô����M�G�D���B]�:��E9V�z��G�=מ��A�9�7����6�[Uyʃ�h�#�v}���\Ŭ�W��I:��� �*�C�<2 h�Y���U����P��Z�1#���7�1��4���-"������n�Q��/���������Xo7f8��I�̕Pk[靣ľ�.*w F�Ɂ9����ҧ��ĕt�T���>��6�W��A
�B�6��YJ��X[��*�(��i��_炥K�+��O �j�tnS���{�bn�_� R�zS0ң��F�
�B}��W��NÉ��vz���za��L*��۳�5�G?��V���[m��?%4�d7G���Z���"�1mze���+u?��˧&��g�T{:U��AF�G����p�\�t�'X�{/�.H-MO���I�O�(%>��mq�9eѳ8�qL�Lخ�(����$��A��`[�F"y Gl1��)�Tyx*{R�2�ތؿ3-c�(=��E7��ZJ�?WE�OF)�鮝:�W��{�=������`2_{G��:�Kɜ_>�p������T��BZ;�</����tX�(�=_�л��9�ݧ $�}� a�r�������Ymռre0�o������U�M�ɕ���ڶ��ꡬ�D˜@~�3�~R� ��ZB�Jc9O/C�:`l=!����� ��67�#���q2���f7��/]+�B�m�%�c�/Xu��I"2�sߗ��Z�����5���>]E��O�N�(���Rx�����xc@�gI4W��d��x/���{�NإĢ�b��o��ak�b�|�h�S���,�����@��^��g�Q���"�f>�}	�^~�A���q�>pH�R�Ɩ?��w�Pc��&�DN�Tft�����W��E�� �ą��?҂[)�S�)XG�I`���\�{g6���=��_
 L:���"Q/���ʊV2���Ft$�����q[8���QsiL�$�]��ue[s2xՊRᝄ��`-���z�>��[�������^j�7W9�=����@�t���j�WI�<��%T�JD7��_��_�d�q�����v�1Ja�R��N�
���r{�p��'����!�F����������V�ؤ1g�k�� �y���|��˾����s��R.5їY2~D����0��P�Ͷ&u��(AR~�N�lO"��
�8�h�����p�������[\�(�0�j�a��|�>evL�̱�����+lFZr'�>�7��@>���Y}~��QCr��&z��1z��Ο��O/��x:z�v���Hb��}ˀ��}E$T)���Q����Eæ�DZ/�
��X���i}QG�E~�,�("tT٬݅�)kc,���K\�.g����O�6�LooYX���E*�St��q�BW�b��z�����D<]hݲ[�M�[�H���w�Qh��U�5R��
7�oVL����|�M�D�{P�t���V�Ȝ �����Kb�ʕg��01X��-$�r!�������I��ꃿ�}��œ)h�V-/�-�`��j�ڧ~��D(��P9��X���Bt�دuٽl���y�()a	j17!�$�w�4Z\8�~����
c�yܖ&�=R�KՐ�'C	s[�FI0��r(�=����T"@��%�v��)�"���Ҟq�
0��l�7�{z���X���}�
sO��MK�ø���S�VE�I� 0Zh.L�GE��ǻo��0��#��� ������Z�AtM5o8<1�_Q����|�k�������櫉t�(�u�P-?������i��d`�����UYu!����n(�崽��<Gb1��Ĝ�s�H�t��ދ��R�kx�^|��^n�h0�����ۦ!@�ge����x��;���Hx�{����Q��������\��K��Y:��.���>�E���j�x�J�c*�����܇6
z�͏b��`5���'��#Um�$Hw�'QJ�x"��`�we~6B4���t�mX&{�MQ�Ȍ��db�P;W;��>���}��ڇ��z}�hS� �C$�w!/W�V��w��]V!C�5|"K��}��Ƿ�T��X<CS� ���(���
���Ϳ��B�_2�/Z���X�� qr�0�2�,S5s�ݔ�i��y"s�7v1��E�*.�)
3+",/Emܣ>G�4o��]���3O,�S�:�����L�iu�!.��x�'1���c�##�!��FE�8�"k��l������Q/GH��~"Փ���"���p����-bLO�2F���KǍue���y@2	8#|�9�3�)�g�i�"�+[u�y��ʄ=��o������p`����El��{��I�qx����Fq�?i@%�'ڞ	�EpД��M���&$���H	G�%��:����w=���F4����_��dW._@}�<k�D;U��A�\qB�9�j��e�e"���B��ã �#��c��F�C���힂 �9(�Kq]]VL��}��-jx�y$�su�aTzAl�����m�-eA��ȀO����4�L aNvWao�wo	�`;�f�y��p\��]<�Vv�1ʀ!"(䪪ҋ����B4�Yѿ��7f)޻�9i��!�/��ot��%A9C`�ѿ��B	
c�̞�s�I:���+bY�U��©��5��FR>�[?�o~���vu0;�[���F\��WGB�vO�����S�Y�!��b<�_�M;q'�$W�fym�@�i����<�bu~@Ğ%�غi
�3{�B? �mA?m�<er�ҷ��E�.�e�*�[����P��}Y��C�n����)�oZ ny������'�z�¼�[醲���/�XG��/M.RW3'�i�z��Zx��t	�74�.��еD�����F3T�,�:�)���5�����?�w?	�9�|e�����Ćy��<�J��C�N����_�A�ʚ���Ouq�U4�&\��_cy���}??���.��
�V�u���X�źC�wz�ڃ8��n]���&�X�y�P���}a�����{�a��])���vD�
���D� �2E���jXsJڋ�%@n�"�E?�a.��xf�[D�����ۣ�`>���j��[e�N��ӂ�W8���u�R^���d7�C���O ��q����p����=\�eu�{��v�"V�w�a�cU$��A�o�ª�'�.ݖk��h'6��vC_5U��AV�b��_�?�Φ��cd��m-E����������L@�%X���BG�����Ô�͌�T�%�T��\�K)(ȮŴ�x�,��9J5�	����,�0�r��N�q������ӪZ��Z�A������}�f(zs��V&Z�[G�l����dUI�v�$�|q]C���ha�8{�*�P��//���]̥������mH܄�{�	�I�ػ(�6{�m�U�}�kfN�;�owao|�=kȕ}����˯_Ѣ���v�7����{�+0H��>lڠ��m���8�s��9S)��A>���%!z�dU��9d�����B[��B&3
%�PLT_�Z��yt�^��7]��6�޶�A�2�%o3�R�����>\
Zd�g�Y,�_j�z����V�b�] �Y�K,�Է�c�>�u\j&��D,q���@�X4C�6�?Ŷ�o�����5~�P��]�w���+����
�@�y�\����8��I/%H����I��]�7�P��.�X�,�G!�F ��������SE72�U�{�K��U������Tg�z}a3�?��d1b_]�@�`ٹj L��u��@���T��.�� 8�K @�Ǿ����+��P� ��瀨�!��u�gl�����V��y�E����Z��<��<�1��<R{����T͆��0��4��ǃ&.ZV.��~V��`ڈT�\�fs����4�`�vVp] �f>�[�¸S����5��ע�����qUC����^Rf���*?�Nu*����򒣖>����ě�t��l�^xk�ߝ���2H���3����2�]̾��4k���~+gX���x�m:�*yR]i��U7
j�5�������c�8#$�X�aаL��'�0| a�2v߳ ��0~�D�?dX��R]��]���M��+�,�'������,ߠK���N�0�s�u��.�e�D�� �4-+l	���
筴F�۳������5 =����O[?~ܦ������u�@%�����e�u�����L�-�t&#��kjj�U����,@��ƄT��P��i -�p�^?��S5+"�q�<��;ׁ�b#g6�T���pE-��7��UT���)�.`z�`t ���$뿨xmJ�ĕ�O��Y^�Y��3 ?�vċzoУ	p�X *$�D.��%=mzVRu��"C��*H�E~��R��:9V( QdK��<(���7>Yp�s�fI����نe��K�پ���ͷ;�Q�<���#���	u��*1�����q20��u&�}K�O5�/;�J�R[���<�+�Wl�`ډ��a���[51d.��g�����#a;|�u��wO�Hf���y,���� � \	K�Xb�Y���/1Ŗ;a����[U�Б�/��Cs��ͧFJ  �߳��7U�:_B���Ɔ�B�G\8!�ѻ��8'�pR ��#sXlxV64EB    fa00    2710k5";s��"6f�7��G�*���l�ؚk�5(��+��7���S6b���[i_5�F�p?S��G*�j��qr�(��f�B��{а�4�S@a�F�"���6z8�`����h�`|P��/�����{������z��$�g�?k�>4_y8�YLN\��vOQrS�̧r�nBBޥ�;rRd���T@�h#J1��Eɽ��V<�J1��w�zV��'v��іU�5�N���?,����pο�&)��ؼUl�KQ�W0��G�EuRt^����@;�t��5��3�� uv�N��k�w(,�� �`!
Tۖ������~zO�&�]���3�z�J�F��_u�\Ea
�@V�d��˟�1&S��W<"��9���_�M����ʑ�5�O;U���KCd��U!�'h:��?߲
��˨��9V����ȺYԩZ��@�S9�TN�.����q!:�.b�m��g��,ϼE$�=2`��/�6��jZ ������|�=�[H���#0/�|y6�.�4�!R�Z���;�g���_�J6��`�;X��۶_�7T�,�i,}��E4f��%��Y�eݤO�J��T���?S9PF^�M�G��N:��df0x�����`x+�T���$sĳwaPB��r9��J�$���T2!ko�^�3�l5����b�7�����M`��� �L;];�d���y��i�D�RqFg�T��s�P���e���yZU
.���S,ȉ��r�b?�[�Hhb�l���{���߾=��{z�\͒.���6б�g U�j�h��.���b�.Z���6����T !U�'d�y�Q�����J;�3l���_^4�NB�'sYY+'f��/b7��¯���B��f���\��8h�~�N����w�ڱ/���lyN~8W:  ���ZJ�T��:�CdھJ�ٞ8�!����t���;\�BG �.�S:�D�֞�C��� G���O����l���ǯWUܨӳ�p`�╄�W0*-�a�z�M��X��p�7o������sP�)ԇT�%l�Ǘ_؀g�)S(_|�(����G}��?�ӱ�bҦ����fg�PAQt�v1�D;'^�����4ڟр��^�;�I��9ϬŎ�+�z��7�ӸC����+WT����)���'8ْ^	�A�v,$��R�P�M�p�^ht�d�-
�/�=�_�΄G���1����u��V��bh]�jF��fOzVq7��*��|�w(,��&V�(�/��*��u�:j�S������s3�U$�$Hk��R���Jҫ
=����:`��nd<���4V8ʴ��ﭹz�JY��a��㑁�;pP��=���������j#3�﬙��su�Ej�q�~,r�6Ꮘ1Ԅw��a��@1�\����r�
�"l�ƕ2��R�(���Ғnđ;v�ߜ� � "p�$˛&e�#
����{A���/W� ٛ���@o�����i�V�t�ݘ�g*�k�Ȼ��)"�@�^rNO��x��B⼓�a)��[�7d�l���������dl� 7�r�р�T��bC&u�1^�'�zR�Y�Ys�Mٱ� �̊��a��bH8_�+|�]e*���Ԣ�3uf�}�}������L7Z�"��`�.l�"��k���.]C��b\A����	.&Bkb��I���F��>�M��(�9�����=�Дa�=���z 9��Q�f:�\/Ɵn��G�g�I��C��Mxnqe�=����wD�{>����bp+8�b�	K������+v��J�s��L�_���v���(E�V��\L��#�sn�j�jYY�L�I.�;)utMBp��VRŲ�w'�X�%}tb�ǰŲ���J��b��C�R������+y"�B�|u#�����|���Ec��T�X�J�/	s�v�Ӵq��^=f+��)�1l5�Pnn&���[|�o��������CˈI��,n�����|�s��+Y�?t�C��;[0�^c*�k?���*σ�/��EV��H��`�aO�i�(ħ@L?�beO�Ɇ�/�fS�����Q��C�Ub�.R�G�7T�&/Ӕ���8�n/���W��r L���i��
�D9�d�i����kg��� F��8�l��S�|���K�Qt�+�#�������m�?̼��PT��EQfZ�|˗UO����k������}HF��OW��9�5:csT���ٖ.E���ѐGc[�MF��2�ﭪ���K(4�QW�(�^��kK�P!j�6�l����Cx�VR����p1�{���~Yo�Kh���Sb�F�ލ�=xõt�q;#f��z��"'��*�Dlwf:}h����g'#QZ���[���zU*8n�����0����L	�R�ܝț�Y��p}�	���0�dv��1$孶�=8:�9��τvd�m�Fq�-9{+�K����q��5�:��W.���u:M�q��Y��	|j[��Gf�å_��(ouB�fq��aE����˳��!�#Ĉ٬᫒F�����%�֬Ip}kM�YWZ�g���E���Q�r2.:�_��&~��Ux��u���FʴO���Ή��l����	=���(r�)��op���64�@�o���,9�I�
�v�5p!W����|���ML���X@@���+��������9��U�(F��;e9�QZ�7tNӡ]���Н[9v5QV���?�96�OO��1��׎�}�H[ۧ�?r�c�@��ܭ�x��r�$�&���nٔ�X[ H���.�r����xi�`Y�϶1�c[7��m��d\uG�K��W�P*n���+�VJ�?V�<c�y�՞z�s>�Keƛ�:�����뒹I�RH�r<U5�����}�D�ivJ7`z���Z3i��0Q �G�^q ���6��t�	 g�������I��D�oH�f=�Pe��&�ay�~���i/�@�WG���1�qf}�.�j=wh��Il��5|i��3��d��CE��#d`��L]�`����xcݽ�5 }�����ki}Flr7�*��V-u��<+��R�&�w�¦:Q~`1��̠uӂX��^N�#�R:h~ ���}#�3z�ʹ�ܲ*�oK,�S�M���鶄�
%s4tr�:�'uӦ�՗�a��ن��n�\�bl�=ږAkk�4��)w�*:׋������4� i��7R�U��LPn��<���X.5�s�y�����Gz`�r���MyI����g����V� �p��,ȫu !#'Ǡ�]������f:���^:�	]�"V��0�.�1&^=r��TG��Z�yM��0+#��w̱2̒㵁�Z�a��H�u4�)���G��@�;'���DK�?31X�D@�i#�ܟ�ވ��a�*c�]%��yj56qG�{�|��f<��T�"�4O�8rlG�8DR�]�e1��OB��H8�rF+dDW=[]?mD�m����XO���tܜ��<���1D84�Y�tx��+���(b�?�78qw����ͽ�ޖAWU�ʅ�$�kkц6
)�Jf��sQ=�UR7�.󈡪 �SE���i�ϔ�@!/|��z��|	�i��:
ߚ$<�r�)l�e}_�����f�^��,	�k��Y)���s��g�/0�����M�x����'^�6�8]�#��������<���B��h������=����br����.�]�%N%`�Y�EC9�m��6.�es���m�-ۍ;������j4�s�:���P>�є��8�$�?��
�ͦK��w�}���FVH��Bg�.��~:$�G}�}50��"ji�Lz����4�J��]P	�k��%R.�:;j�y���Ϭk�F-�NX��C�(�ׁ�2�Y�N>IR�=��_Cܷ����7�}����Hn��z���+;�e\�?U�����+)��b�S5X��HFn��R~�7�w��T�&����f��Ih�F�g�����MZ��W�x
¡M2e*���P�)F%MCz����sG�t5ykj�E^��f�NB9$�Zh���NT���qNv��
����JWٌ�9y�g��_����ͤ=J�ţP(HF��[p��h��E�� ����i�cܐ��t��-Z\پ�Zh5!I�t�U��7�,�Ѹ_ʠr�zv����6s<r�+X�#���R��.w��hwCg{e�W
Й��ԏ���;��ټ��8B6�#ɨ�=˶5�֘h��V>�$�b����Z��"D�WK{����z�5:uEU��r���]q�^�Lxs(�Z��7ts}]�9��~i)� k2ɨ��7@gh<�MhZ�H;\�OrX����tQo���!p�aF>r:�S��9x8h�}�{��#���>/��TҌ��6 �R�>38� >��.��Q�\�I�� �vW8;�C�����U%9�D�p�w3��=jZ�i,��z�~'��!^Vɔ��vM� 6�������0�e7��ѷ�����Υΰ��_��h���ͣ�/�$&�l������4�d{�1
 ���πĘhy	/@�(�R�c4�� $��ߍ�E��/�o��x�Dl��������V�X�j]�<#ɦ��_1�Ґ�,*�� k��Vp��*��=A^!o�ͺM���4�N�8��"!�y�0jU�p�5y����+j�����s>}�
#,o�EF*w�ѓO��:M?n?�x�,Ft[G����*�v��KO�	� �OGRC��Hz eu����'���e�_X��Ӑz�,����x�:|�,8,��HP��",�Tj�>�&D�=�!q��,-OjF���<�F%����(:.Z��!����rcm3� D<���H���>�D��lDh���T�2�H�`�Ms�St�䂩��؈\@��>���o[[�E�JX�&���E��o?�M��� ����C!��`� 3.u� �t
�3�� ��c����������rt�>o��[@�wץUea�jn}�3��^b�R
���p�8��f�+O{�7�o��p��35*=}�R��Z�>`��tQ��k�$c����NMZ9��h�ވ%q��I���g��/e_��-�N%��&�C���p}Rs���)��:}1�/�:�7�+H���#�JZr��pjS��|��	G�g�L��N����*?��� �y�d�K�Z�a��9(���Y��9���Ɛ�
aG5fL�1�̸Ԕ��R�<͗����k�Dl E'@�1��ak1��--�3-�%�^�U�ERF��Q���m�8���xo�:M<��ʤ��_�pF{�b؃C;�`ٸ?<^��p��cB c�'2DJƦ� ��!���(�~��E�z�(*F~�Ӂ�rS�j̘y��s_,�Y�F�
ҁT�s�W��}�Ћ�<������o��/g��n��G������V�}�u�/�d�4C���M��C�̧[w�^	�r!�Zst�I�3���Qs����ק&��jR�p� ���a���m[.�jI�5 *�Ԡ�C���HN�>ӂ~�<f �I�ء�>%	YG"|�}�ף~���f���@�.X0Soȶ]o�����ue6_�C�,�$���΄�����b�k��9݂D^��ݓ�����Q��!Q�!���Yq��_B<z�#b1��3��k%�����h�lBj.ɚ�@.�����`��ir԰��J��e}"w9�v%�8P�1�Gge��Ze��H��>@�0�ջTвϲ��0����=)�G��/w}����gW^��s����_�
�xȶ>o�/Gx/p�l��'P	su��3��,��u�v6���\� F�K�Z��Q�CO�H޺F�|��-&d�����k�?7\$�-7�t>'���e�Ͼ�����Z7��rC���phq���9��X�v���yU���)��L���-|vu~�H�t�V��ݐ�� ���Yyn�Jf|Y��T�~�0#�JL��yU�C:�-_(�˪yax����\7�P����:��|3"HF}�Z	��}+�d����~/+��[�6���v�W��M�#o"&��>��Re��A�6n@gIJŞ�3v�V����c��D:���}#��]Χ^ŕe-��)gR�gc�]�WɖxCwh���Y��_Kܲ�ZEʢ�:�2n��T�I_s�Ԙ� ݒ���'�@��}i?���a�c������%ҝ38�Yuf�l���tnX�*�Y(��oh���o�v	}�C��o9�Q6�J2`�y�]`ݡ
�to~I�[�K,�Y�=�5�+y�ߩ*=%Lp��	?�-��'��Z��FWb��EV�,�
�����A���9��?��ᶒ+�ӛ��H��<x�o�F�6��V�F�8�\�c����G��O�h��fC��/��}��+�s�v_}?�����J�10K��^i�y���)��p�E^��OMUat�-��n�K��l��Z�o̢�i�(�*d
�x�է�Zۿ͓��6���Ġ9a6Dr"�V!g"ֹ<������X�����@��=ĸ߶4�T{ꡏ�0a��^��E��q>��<oE���]�<��Cj��`�[_x������w�_��n�xf��g�p�n��1�a�>ɉ.Kh�6������E+ G�3���@�3A*�N�`R��u���D���Y2U�4!��Ũ�E��;M�i�jK�&%��8��o����/0���Q�X���$�b ��c"��m�I���ʂ�f����1m�`����G�5�oH\M��U�h3J�8X¹6�-Z7�p&�})�\W���U�c�ڢ��9tf� 4���gkE?j$՝�OLJ�.�K�Rj-�+��h�S0��Ub�_9����ԏ�W��Y�Y��#�q�V�y�4GA֩�ѹ�g�����+�I_�輪��{����8��=�\3��JK;���S(AS���)�p��}�@R�հ�L�S��m*��W����5��=�s�����6�blߚV��˿Mf[9IH!������D�eW��E#�<�^G��
E���tS��?vǚe��-��}�!���7j�)��2�IU���%�qhw�jU{�0yYڳ��i�z���}1�uf�*�@Z�s�,�n�}�$�;��2D%Q3�
E�Is��5\K�ۨY:.�?N�1w����e�t�n�ʜ![�T�=�eMGp�yQ=��G�W��*�4�N���?ц�)9v"8zD�POG<`�4C%�������Z���SMY�3t��Q�U�C3p}M���8h��6B/CwN�kuƱ�С�ZdQU
RܠF�]��u�Ƿ�&Q$ݱw�*4�m���t����Ë����G����A�����8�Q��w�|����C(Zl��b�����R� �Ф��xS�sC��P�"��o�Oe6���^1=�JD�%��C�����(�VZ��ph��8C ��8k;��߭�E�w�q��/&bw&)nҜ|��\z�4e#{�(�)Z�F���w|Sc�m��l<>*�! �����;�V��b�uQ������:����
��3�o��_���V�:�\|��5]������_T�^�+ӓ����
�z�����9�_�^|8�v�V\�iO'���f�-���W�pz�
E��x4%g�{���P9.�ʒ\/0ǖd� G�3\�Ԅ��0�qO`·
���e�=�7��,@���C����Z`t0/x�ۉ�z�=|mY�D�®&H_8[>�Ef�)F�_��$�V�H+ᗠ�q0�y�������0�E^��Y�l�RҶ�����\�#�.��%��ȉ����{0��pc[W�9wk0Q��p�t�XI�X�I�JCػf� �[J�Қ� `�����H���-��
}�?�j��.�,!|֩"TM�ċɬ��
�ۛ�U�� e��q�(�uJ�;$��\e冞�9��r���Mb�tF��a*:�_����C�JM����M�wB�&����s�x3��\�s�ޖ7�5�oAa:�DI��'�p�Y�>��
d�� �u����xLl�C��
��1���N�yt�F�e��R��j�a��akh[Y�\�G[?�e�
^���t.����65�M,��58��T�"�??�JDAMH	�P��'e@�TKłN�q/��]�9�~���S�9ҫ��\���ԟ�T�f���>rt�e+��Y��<'������ś�s
�7>�V�vO��"|���rxJ��Q_��B!hʘ�a.��Ĝi�;gM�wQ�0?}^ˈ~gx�t)��R�a�M���3�nq~P{@폘g�oG�!s_߫MMή3|������)Wyj<��> U6c�qD�����Ɩ��z�����l�v��~�n?C�'��;��*����E>��)8�����H�r��Q�\\e<j8uɶ���iZ0��C��$�K�:R��i]�%	���=��6��g��[j��$��@���	�����$/<#�{�(�"�A��-q��?T9����+O��B��n��f�O$�7���3�����s�Fl� ;4�e)�����z���ў�╝�x�+* �v>���/�#+>Dv;��$���S}�7��?��0�+����1W�2�O y��[ؒ�$ڟ+Ehg�y�
�啤kw�����/IY��������0uD�!l� ��ݣUn�˙9�>^S���~����͎}�3�f�Du휾yA	���f�*��2AWg�|vh60�hs�x��O��h�Nk����.n�Z�=���;��TS��Y�f���3,�[Oe�	ᬚ(��G'��j��ǅ�7����G06dD*����20LD1��a�ƍQ`5����F��(�Jp6E�%�?�,/<e1no��P������
&-&U������=�zn�J�����zʴ����ظ����x=vԵ���u����PhQ�2l=�=��/�uH��퉤gF0��ңۛE
��WԮ�y��4��	��m��6$y�k��ڲZ�{z^��G,!���i�"L��դH�A�XIHfd?�JJ{�q����b�F|c�:j��x쒢�����ږ2��X��*#M�:z��)ƦQ����T��K����� ��$u����"�X*���N"HX��`Bw�%j�L`��sp�3���gEH����b&@�����<�me����R[��<��?`�2���z;�t��q����+%�w�O�sP��^E�?���AC��K�h4��������T/�jQ�*�yG�}�c�s�l�S@�8��s��P
��R߃�|�л�ϕ�'ܭ�zk�eݐ݊p]m�zT�X�¸�����M;��)��(��"w�
��աJN�k�2���?��K��e�������W%���bwk�#5���~����G11�f�֬����^�r'�5%!@u�U�|ga�1�7nF)�13��5��+��"��/م��F��3�%�%�紲���X/6h�o_��a�Ԃ�{I�����'Ȗ�� tW��{���t��2��y�g�[v߾ו�'6^@��V�/�&�^��|�6���F�1��lP�z,��.�tn�A�� % �~[�'��ۓ�>�g�.��d���yD�F��ʁDWKЗ0��G��"zt�,��yLe-�VG��π-�c���B�4��"�)x
ReQ���[�Yk�yi�O�##]S�-ɹ��ONF�����xZ1	�"#o&c����:���A�tA�[c-'~��õ�K�Q�c�dgh]�o��陵E�v�=���\!����J�����R!1��g�d��'�s�h�&�q�KQ%|�/����였8hu66#F6b�?#'X,B����>��_�pZ��~��`H�d?[:	S2�A�|�Y={XlxV64EB    fa00    2420�'�p:�x�i�?~�<��^�Z`�1'w�K�^���c'��P�+�ϾFH�%�!�(z�����׌�ǣ+}pw����Ө�vӊw�a���������W������Br�Q�z����T{u��N�B�Ic2��>X�ZU���?�����!���M4�J��`f%�� � r�W���|����:��b��Jա�ɘ]m-�	G���c�D��qW�f�f1�Ö�Q2&���w*��$�X�J7��hs�.*��?��)m�ÍmT�&溏%��
�b�x�CP%J��U �l0Z}��?A�u+�	**��ҝ�����@U���\��P�O��1Gη�#rF�/3W2���:{�/�j�)FO�P�ܪݾ8��$�܉��$ߏ+���dH�Ԭ��kH�Mm�0��BRIsѡ���+!����✕�k� a.��7�]�3���Y����{��g��{�dDI��%����+����]��A����������h)%�G<u*Ⱥ�5��G���D�Ǧl�_j�.�2C�?�ZXJ�j@���� �bX�=���'PȺ����@ֵ�_MՁ�R�S |�v��y �}�DV_�1nghӿO#������-�����O��1!�ԓ0 �(��
m��l,g6˸r�ov?yО������P�6@��O���q�1SV�i�Ol��G:�Ơ���9�gks�Y"]̅��.Y�KFʨv�
w[��Z���F.M+�M��ϸ�xNA�Jd��$�1��3�[.�&�0�Ӱ�"Zn���������]*P��'䜈�:�Ϧ�ݏ�;����Ʒ���))T.G�ʁ
\�4Z�)�NC�wo���qk��ts��q���]CV!�d{��u��щ��ؤN�΢#.�R^��m~R�Qt�a63i�/���'tń~ޘ��`A�T�Qa�c��s*C�����\ƞ'֦�"U�n��۱�(�dqgq���n�K�g�Ń�ٞ��7#���.|x"u�+ؙ�im����&\}�uQ["�ͦK���u�]QG���y�'�Ui�~��T�d���Z-�Ͱ��9�\��&���������ݗ�1��Ϧ� ���a����1V>B7��}�û�w���=%ǟ�ݲ)4��� �#6 �b��&���<��+r[Q�rR��!�/�Gw]�̶h�_\�"�{�D�`~�|����;�=�=�� U���}�y�[cd"V�NO�r���� �-?Խ2Z�Q|�_��5���b~-�\���Z����$I_��[ �;L��ʠ(,I����X@@BZA�����X�a�0.8�����,y�ʂc��2���'*�9����ϠH��nCT�*��M��;�1Ƞ�v{���&MyuP�՚����9��2�l[����>A�czL�4�����$��*��7r�˷@�|\E���0® 
��ˑ�+��R�~�.d�BC�Y�Q\�=�`���*έ��{¸v��{�"M��lI�	&Ȧ���A��FgzͱTƇj�4�pQ������G#��M��(�`��������RX�����&�cEG!u�����mԔ瀇�̀�,-�5�f���(x��K�`��[@�=7t��,.Ѻy� ��;�/�,
��Mx����Z�l�;���H8)��Ί��e|�D�{z�dg3%�,A`�g�TZ�5_"� R����0���V���>��򱮉��8o~������w0G4��y���享A�{�AL��pN�ޛ�	��
=���ƶ8�r�*a�VG��ly�E+'pj޴o5�;��2tQ֔����G�'e��yY��sf9m�P�#C���mm���D�}[�*�H��O�:��PO���+��t�M ID��$�6��V��a�9���M�<
�M��C���L�|�����b�^�x7iJ�P�sqɝ� j�C�ܩk���Ω�˱�g�}�MJd:����� %M'�X���*��~}��Q[)��W���,�0�y�x��g�O�/<o����9�2��4����(�J�_gr rå�;ٶ������Q��7 \�*���腱ھ����%��Q��ԁ_��X����ܡM�De��t'���-)F)�g���aLb����+!�=�����r��k���8�R�@���%����!��
^����:�I�&��kI�O� �KE��R9́��������D�:��!�f�ƆQU�]�w�&7���#�>لr��<6�!����3z�*�-
p2	e���$&NWNQ�e����J�{R�W����F����?/���V�(���˼Lw�Aw9".V2�$-ܶ>�>��R�Pg�1���h�6�\x[���y)��mZ����h��J;t�ڣ�*��S5�Ȝ�ub-��h*����M+��+n�&����{q*�N�9f&Px��ۢ�8�}F��BAu˂��?�z���)O�%�5��ϊ���:��Thxg}��:�KLfXTrq�%�n���_b��c�=��ig�5SzΣO�6��_n��?���l��Z�����}���v^�%g3^�ǯɸ�l%.ϒ�6A+α<2�M��mo��N�&�w� �J��ml�i3���0���n�:�bm�e$��9�$�cO��}չ�:虓�!ٟ�pz�d͓�mmwm���l���� ��y�����&��0n���bx�W@�[
]�>�����8Ľj{�잢�g�Q%��2*:-�����x�+�8� �^�>x#��d���a���j���,gx��i�?0�aS�~n���W0(3��h*��xֳ^�C�^���S	Mt@�^���7��~����]X�M� �]nO}�	|A�	'\�ȗ�Ժ����o��X��ˎ��r����x/jT>(�g�8�����C[1�m�>������Z����_P11�%���u�
�&��
���'E����g�1��E�Ж�^b{�<��&��C1)a�K�lʶ�ܠ3��*˳����UʿyǮ�^�%�V��:����&	���˞6.��
�ڠ SM;�����z�[>9���ےc*|5!R�'�|$a�`����9���N�����;�ʶؗ�ӽ��>�!�:7�z�%�F|M�y�����a������N�����i��7ЄPj�=�%�=���]V�Dߝ�Y�#�wZD�$��<���Fz��
��As	e�Vy��r>"{���S��<�*�� �
h�4h`J~3e-]5��{Sm�׈�R����l�BFI��"\�qa�3z���A�\�W8[84!��b��&�Y���8�9��ݯ5�/��9o���YO� '��Ne���Ԟu���p�k��y�0�ں=��$����ÁXrCA�S��8H8 l˭>S�D�%�u��9��?���
Q>OR�^���C��+�Ӥ�4��\B�m��cfτmџ�-��HxbQ�І�]|��"�.n�2s�g��}qD���8�E�w_��LB�ų:ͅ~��Ms��C�Z`����J[0�j�v�������!�6��X+��XM>��_"���2����"�N+�g�%�� ��Z���:w��������OP�V���_$���t�&��!^/}��od���P2�^o��5A��=T
��I��|��j6��_�3k��[�ݯӌ>�>����_)��J���T��aE�3�heSob'�s�lK��RP��8��+nV�)�.�=�b��7|+E�Z��oJ��V��	�6Ҭ����rc�
��`L�ץ���V3I��-U� V�[b���c�"9���q�:h�Z %�0ݕ����{%{;�{]Nަ�i�)�iR�=?U�gO�i�����j�&�r�R��y�tV��e �n��Bd`���X�F�#�����Pl)g/��R��Z�@������i��U�G�h��͎WCZa2[E�D�VZ���� Z����ʐ.c܈ ���~h_�'���̥��8�:��	��郕}'eC@�����������������CF�F�=;
�)�G��@i#�:�B�27�s$����ᦒ�2��,׃�X���pf
~�`�����5ހ�|�*�<d4���>4��NW�O9Z�?�w{Q����
���ئI���<�=ξ��>��|�>h�'���}���]x����d�֎����P���ӹ��"� �v�vʞ�-c���2$���%�v�$R"z"2��}����bp��RmXQVA=&����~W'ѤQ�"��%���5��0�[}XU���Ɉ3����J�8�RfK9<�w��p����V��z�|���>���pW���4�6�`�ek��# ��ɲ�$4�9�S�
w�P�(T"�K���tA ;LWU���ª
k��%+���|�l�& OXՕ��?Dڃ3E%������D����Q��ٶ��F,�~�<	��-\N�x3�ʯ*�3�aIC�[r�}Pr̻����Cv�n�߷��^�5��_Z���K�a�Z�դ�Z�
�4��(0�>=ǹ�����H�w,��z��[��(溮�(���>���r4�*��!����:5����x�aI��5�e���$�gV�z��ټ��Xu�d��4_+Badͤt;?N�zL�8�m&�P;#8�u�A����G�:�����~4���m�rqa�J��.��CF/�����Q�����ӝ���M�b0E�$��Eg�F?�`X{�J�GfN�vtT'AJ�w�>#�� ��.Jd��V� Ҽ��L�:��)i`މ�#}�Y�JP>Ǥ������]�6��Nm{�޶_�RġJ��9P{LRn�����6:��.��;�R:�i��(wBwEԟ���>r@������+��j~���`��W`���.�a	W�e��S��O��@U���)5�z�=oTā�R�¿G~H��E$��C����ǎ1ە�$DM���}�e��Y��P `�u�R%M2#8��'����ܚqo�P�K+S�pOQ�(;�Dr;�@~[ӧ0�i�<9a�W�_�?W��7�[�|&��,<�t`�v���(�V����y��O�ؤ��o�S��;�KƏ����*ZXDfČ������MN���Q
��ꭥX�"��L�$&�$=��`M{v�{�L+�h����r�y�]��i������"�����9��̈�ec��]uٰ����Q��zM��$�Q��l����s�#����XF�IW�?�,Yh�[�}�I�{���<�z���*(���7Gp�W@�1t���>��"EM��L����P?��-�1֡ŉ��bx���2Dù�ʞeժm�H�k[*7��u��7X���K)�uyA��`a���4#�i����
�h��TJ}��}iR�Tj�l�%�H���Y�<�Vt��2��(L튦�������Uq�v�����e;u1�Cӓ8c>K@�������.h�����9O���ȅI���TfyY�q���!�x��!C�����X�*Zi�T�D2@�Dkr�:��SV|�ɾ�;��M�,9gX�G����fy���4����_��>�h)�
�_�����ٗ���
ex����S�h�G��KNݳ��eyC�i4��Ak^�O�v�G�(N�󴙦���p Ʀ��z����|[-
Wg7�f-P�sQ y�-�2�ץ��c+
��ǅ�9�e��5\ �A�eݼ�c �-_�-�U�+����?����-��FM'���iġw�@��6�߄���\ ��RLZփ02�ռ�9�W�N.���Fbw]u�sz�`��e9�v�!��{��a+z��{60���|6%�l��C���'�ЎM����=��)�[5�Կ�j'N�����t �!��?#̲x�u�>�HdQz]0\Y��b�7���!GP��6R�	�N'�\�E�=�0�����i�1@7 �N�im�G9ҽP�I�	�0�˦�T�ӋE����LЎ�1�k�!��_�%jБ���89�&#��f�T�4,�cVYD L��}��1��1�s�K��e�Uf��؂�����ڡv�p��|�r�����Z�vE�$��v���x���Y���#�P���i��S��D���m'Ŝ�>�OM�P��@ �h�A8��q�MJB-O^���cp�cf�
��ӌgC|�� а�}��J���x��	"��8���JC2��D".���.�
����C��p)��!�E�8�®N��'4�h��_WN�!$V����2�(t��V 2K��1��&����cI�@q%�%
Z$��i�bf��c�+����E��i!)۱���,
3/���#�v8{?���'A��`�H�F�D�gv�+��^	2Bݕ�ۤ��=��]����p��гB�	�{��*w�E�{��~�A���t�0d��C��3A07���H�M�b�q��Sd�,j�+s���ҋ)竪Rv�����Ƽw�JTf�K����v�v�?vᥖ3Wy�z�%���Fw��vd6������Dٰ�NyH3�m�ߒ�#�N����	��Q�MBr�5eCQ�~�Y�
����`���x�Ԯ�R�o��H�!L�`�ψ���]�>�E�>4D|]~��w�a�ps��оkSp�2n�}��cQ2J�m���k��g8.�ho��p�����̒����n��B�pϳ|��)f�W����h�i>u|,ju �:Olߑ�A fQ�d�J8ń@ ���u�����ӧH��� ��^ >�>@T�r�X_c�S���ش�0Bq�a��"}�V�q��L�$�dsϏ�/�-~sH��0�9��++���]�u��c�Ԗ���p�,�<sP��5_�dË@�����ܺ=�rl!D	sXA�s���S��6��e)'��K[ɉ��^15U�欧p�6�:�#�{�<��K�'���7Q�(�j$�I�v�<vӒ�&�T5�'�w�/GKMΎ��L���/��CP�i�d4h.Zgnë*��2�+��fxאLIr1㚗��F�bQ���r9l�V�G�,����ä4�!��Վ�'��f�T˙-��,��A�oF�tc��=�P�V9x3�����B.<�� �Zi�����o������ALs(���||��Z��Ѭ�)�2~�i��@n�f��c�2욹�X��c�և�M�⃣d��%�vۇ�&x�H}���]zaBk½.0~!��н��N~ئW䩚��,_���ɏ_�:r��^u� �7�|d9�Z�Yݡ�Iߓ�DGC����/G���z�#�y��<����R� �9�Gk�b@s?O��v�J9,�W!U��Z<���0	��P�-Ŏ5I����n��Kk_�M�'�}Md�iԭ�{߁�@5'A0��_���)N>,��5�� X�r4D7�Ȉ���v�_��vٌ�as�_A�g�;��A~8��ҟٛ6n�� �z���Li�N��*g�e�_��μ���2���󵑵���Dߏ1�l��PjZz�Q��9R���2w&@��I�S5`ݚ�4.������g�7O��&�g"����*���](��0s���K�j1m�_�t�Abl�|lH�~����j�V��Q��=��H��9{I��n�$��O�DI�&�X2����q
0ͅVNg����ªMY̆�ԹGvAFgަy��?aҢ���ݓp8+�n�]�p'l�p��@�k�'�*t�P���=FZ��g���غ��^��Є��_5�v�Ny�/rQ�@�N�7����i�H��f�nÝ��H�u�!J����0���O�[�������߹寂hE_�`�@���L%�3����ʻ�$h�Eo���UM���0�\3�l��{����Km.�[�!bᒜI���k/�y�c��DZ���Xa��"��n�KXr\ȶ1g��־IְQ�oo��[�M����Jh+�82�i%�۸�HR�L��)]:�0��vk��a�	 ՖFx?O��B3v%�~B��Cj�ATw��0��a��p���%s�<[=��07> ��B,�E~�`�_=���	w?�*p?���.yj~wwl$4.3��8,�c�>�EI#�x���XgF'����> Ѻ���_;���^7�S�bA�����@u�Gs��\ӕ<����1`�sk�r(���K�!��~�w@�� �W��a"b܀ؿ��cx�d��[��?�� �=k�#7.�11�}��i����<�o�� >ǛQ�\"��=^���U�}��E�>�m��5�X�� Yܒ���Pm�6�1{`s݋���8E��m���;��5d}n�t��K���4o�����K�U�%�5}:��q����Ge]������8��L=�X��sDO-{2�<��9o��L��MJ�+�k�B-���&�"<��U�%.u�B�r }v)�$K	�?'�O-��^k:=ں�	1�1y�ċT��k�z\�a���-T~:�x�6�w
?3��������?����������հ��Y���I�v�Y?H[6�"w����dG�vӨ8�j���u+��^"ܽ�Л��fS�b�}Y�\quWo#a��~jq�������L�j���j	#g�[�-����Kg�17�}�n�Ys����<����Î}ED�F���Q0��?X�R!�IJ��pc���wڳ���|�ŕ���w���<#*����6�����=M�h?����R��L퇠�� ��|�i�H½����\��	I�0�>��ZO͹Y+ �zb)Aˤ�(�t��(�t�H�U�Kq����M� "a��Ve]̖��F�?�חQ��i|2�w��t'�ѡ�� 4j�����#�%R��I��x��2�5 {Q�nUΒ�<c��?�Xc� �M����Yt|�
����j������/	)�ι�h�,�<T�ښ�xܟ�F�~�����TC= �5���7ݥ�tBR�5vg��(fC��C�am	�<q�J�N!t�� 3�y�D��DTޠ��&���< ��&��D�-gZ�(Ƒ�Y<����{#9X��iH�ܿ��C��.V�p-�@_h�-@@��z��q@��V��E�@�"P/6 n೒�G���Zv��psK�K���x�/n�JV�1��gg��l�QH�'� ���m}��c���\��ѭ~E��aW(~�}zf�h/���]*��XlxV64EB    379c     a80ޱklKy��L~g(�x���f%:������� ��]%#2�z�!A�^g���A�5�]�������FG
��pq�l"��<���c7�}|#�1�Z]p#�A�C��Dc}�I��r��BԹF�|g��f��s�VEV��6�у�d��4����	�@�Z�s&���,��19����%��������W����#��͸|l}8��+8"�U{�y���=DeF��u��V�ԹM��]�T��rW�H5`pd��kӕ�nl�Z%E����-r��j7�W;���1�d�wi)��	+T���+�� 9VV�v͝�Pk��������� E�w �F��ֿ ʵD�\��r���u�o�	���?�����+(���g���o���h2��*%^��jT�̈́�R�*�n�q^�BOd��+�C']G��������!E�/�5��	��uꍷ�N�\�5Q�Fˠ{��/3�6���˭�#v?�¡�!=h�Z���t#G�A�$����/j02�R�
Laj���Mի�9p��'��mF��p���jŹ�ixe��ɖ�9W2����荔!�?�WؒH����vhfR��O{�~�k> /c�[Eq�%h�F���=����d����>�f���g�$D-&���:�]�6�/_[H�}61� �J����̓�#q�~����Z�@��ۿ(�����0�[�����:��h���4�[3�bsR���c*̖��K$��c;�&>\dY�`��ߠ�`���nd��0���iә
���^<S3���S��b�\Һl$U�J�y�RV��\tV^D��
���`��8��:S�Ȱ���^�U��O��	[�"q���hA�ex�����d�1�J�_�B츝�%�৐�w�Ӯ�,�nI���&��^PLf����}�VN$��ȋ/hV-)S�c�,�)����c	�m����8W���e��k�X�Ir��e;���4Jł�J��o��1�b� �l�xW�uu�	����_�}'�)@�O�?{�95m���,No#{�~�yơ��Θ��"n7�+���(I�x,B-���~X�9�~.a|қ�K1,��/����aƭ�� �y^_^��(֛&��/�߫9��3t�NiR�$���sY�^�e�1#��#�	����b��������|/�� A%����F�s���7a[��$3���b)X�4b�߮!�^�%M���+5�.�et$�Q����d�l�Ǖ�� p�<��'#�1���>��r�bV T��OM�F?6�q������:�YV帆u���r,�0�|��.�ЄP=�8UHx�w��*�[<�r����c���+�Y�V>�ء�o���1�""�f�(\�q��(�����}r�s-u����u�^�Lx�����his���a ��t�����K�����K��k�b��
Pn�K��F.)˨Jd�K�G4Su�1�o�b��_2�u2���m�҅" [�zE(���?qȱс�=_E��^wM峋�Z��CemG�����2�w��Ɋ?2�yN&�&��	�e$K�B�*8�J?�m VK�I�?Q!+k��$�G!9`Ik"�jpaqg!q���k/�1	��k�<)]�\�U�fM���!��L�p�*0;�N��|鍿d�xsPuTn�20&�UUe��t��댲�	�Bm5M8����oO1l�y���o�__�E!�E�-�5ho������l?+�#^�с�1��#:� `��-�"�S���{����G� �\��Ͱoz��#Xʳ�p*���)�53wjS&Dsl�.p���,�f$	��=Q�vx�s�u���������N���r9k���A�.��%N������\��akF<��ؿ-��m�p�b���f!} ���̇�-aU���́Pe���K['R��Cn֪i�$��K��Ծjk�馽�X/��2��Н��#�L�ɋ�.]*�m�㱉NA)�p7��y������(~���%@��yV/�~)���k�<�����8�?ta.%��p�i�NX$a�8�i��?~)�.��b=a�i�c�5}Xg\��ZD�[.�@A���r�u�ߵ�+�rr!��ʗʒ&s_�|5?'�p(�<Cw�0K��,TiG�x�.���c���������Z��_�z�UN��kjW��<�ZX�?♠�h�K�x��Ngp��N��L�}&������)#��C��{��d��)��+����Xũ���+g�)�U��Ld��zy��#=������Z#�XV��9n���-��O��|F$q����\�������圀���I��"s��8t,�����^���;�M�g�K��=a��.��a�*w(� �v�nˊ��`��	3��]dۅ�s,�a#�R#B���p02�$9�RZ�AH�r���m�ñ|��B��p�@�O� ���%1����u!rQ��9�ݞn�Z��B�qo�><�L�L��ϾY�=@[Y{.�/٢3� ��O������C���q��$C���E+縦.��Z��,n;�a��e҇�ws��4�䵑�GV����D�io���1�����X�z�^��\n��������/�7�+��$�vJ`p#���k�8N���E���/z��7h8u�7��d�=������e\VD۰Jf����