XlxV64EB    45f7    1160['��p�YϠ���'`���$�
't��.q����rU�s?�
Zv�>
�CZ�Z������
�uS;Ý��_�	�dHf���*�Mq�^�b><2%�
�H��3yP���%h��p��ÛK*X���-P�Y�Z��E�jͭ�m�![ʶ�kz�
���ÚUY
���rĥ}��p�R.t^7��"�"O	Ɵ��.���-�Z����g���]�Q"�*�y�����L�,#�o�Å�/��jO������Ȼ.˗y&w�H #/[��������8[�\���IH��
�oh�K������-@p�*Z����`�l���:E���j�2l���I37��ږQ��V���F+��ۗ+aN��H��EQs�Rϝs�i��o��h���0�%�^�%��Q �p�c�s6���
4�~���ڴ��)���zRq��N����4��b3�y$���Ui	B���tq���� �(�_�ܺQsH}�G��Zhk�.1�\󐓲��/qƖ����Q�Xʂ`���B6l欥�����І���9�BC_�	+�?����|wQL���*�-G��q���5`��8��A�H.$��{����Ur�F��{Z4���~w8Y,���	{�BG��bS�	�8�hߝM�>YX*����/�S6�>�J���rFi��%t_jv
b���_t���H��b�� ��?�s���qn����vvy���'�h�u��ؔ�uه���/ͬ���O��`y�ur�HH﹩���P�%�R��(��pJ҉��ëӟa���"QB+��ŕ�#N��&�7������I��f'����.-��rj�feJ�b+4"���~ڤNE�|x}Swܸ�n�i��vd��<�?�U��OuV�����,�=MN�6��J��K�K
�V4g��|� �1n�ni��E�o��o7�,4�w'�{��L����a�\E�f
���a
���q�(���H�k�ĺ��%�r���G��Y����m�.'�͢�2A�o3���󭗏�y�ҝ�F�c+�r�\�����e��xN�Ku��p�3ǆ��9��3���{�A�����lӽ�zdWܨ��ѷ�P+@�[ͻ9.I�D{������ ��e
T�z��FU�6K.'�l���'����PqS!fˡ�IP�{j�γ.����%ڟ?C-��d����]:d)���*�����J�S�,�K%M��}�BTS(C�}�������q�i>��{n��9I~�*�!d��fJ�=�J=���T,	Z� XAZ��v�>Mƺ�Ӣ;p��=�#�(�ֲ(4Q;M?�\��5�c<]l���]b���[դ'"���P�G����^��v�f]R�����J����=}��G�+m\��4��|o��*M$@��I5�YGHY*�v�=��Uq�reBח��fJ�=AG5����G�(\f�ʐ�29Jխ�y���E��Z|xa@��b�7ޫت�z�zK�p��c(�nk�4���Zh�+aR���u�hs��*ר��a�11���)���3Zt�׾˞3O�'N��΀prw �N�����F��1�m�5b)in��e�/ludr�����/p��I�20���ھ��r�ê�R���l����)���`b�Bs���\k�����,h��v�k;��	]�����}��M����<�{-�ˋu�TO��&`#Yӯl�Ua;�[,�c˸����'��4�H�V
8>Dڙ�('u�U���$_@����\5J�&s�!��L#P�|���wYk��{vw���;A3�m���&��iaZ��W?2�J\��(Pi��q�7�T4����C,f�P�?B�ja��F4��g�6"���%R&M��~�����w����&F���)[�}��9�d����C�[���H�կz���-�k^r1�{����.sd��=ۜ��E	�j�����3~b��^w�1;�&aؓI��Sm�w�6]�Iw
��~���8"����:|��#�Y�C{��<�!g�Q^�|.w�7��wP�P�9о}�R��Y�~2Õ��;�Z9c�m�<s�p��O|�&&j3���=����T�z�]�~o��\H���C����:��I����~E�%Ƌ��٭R;!yDn��z!�NF����;o:�ܕH!j!7
�v��;_�56E��,��T� �t!?��g�V�p�L��LT.nD����D�l3���ׂVY���^�G�6ų���c�{�C1���j��i����b>�O�s��x;F�l��x�M���=��J��5���������d�_�E��+��,�&���<�w(�I�a�i��Mͳ ����q�B��O���U��+���w�U���Ph���{޻ ��:�$8��B>s���+�A��%�M��X]zX���#�M<# MՎ����//!�s*(3�a�������^ͩӐ��F�~j��JrN��d� ڋ6�6�uR�G�+��Dbǹ�PaôJ�?�`FF%"�r�-Q�:,߼����	$i�<SiI��F�CnO��`�<V sV��@��+��x9�6*L�  Y;���s�.B<��"�s�X�IQK�
��S_+�~��IoP���!h�y)X�t�ef}t#rN�<�a��"���s�B��"k16�ȉ0�C�� �8�Yc'��@���E���❔>-&�#AM���\�	M������}�14���̳u�����Zf}�R)<]1�nHy��4}Ւ�
c��G*��7+y�T��y��V����k{Vɤm]���"öd���r8P� ��}�,Y]�y�l�坣����xI�L'��w�'eYV�Ke s U9z��@��v��R3��gd�����Gp2��Ɉu&
�a)78���!F��m���)D?G ��U�U3���$'�gF��0}TsH�������@�����I�.�Ԍ�(����.ThS��.�μ���;�ԫ�����V/0��<�h�5�]�N��ݔh�*N��˵$���Ucx.@Bw\��D=I2�ջ���n�!(����(�3�R�h��=���@�@���$���B�Ϟ	��3D^��G�V�T�M�������Nj&��Z3̍K��y��'��NT�w�6�w������}�����}[W���q��1���=�t�`D �<�[�������~�Ȏ��w�;8�����HӘ��d4Ҥ��If(6]������@S�4L�[�H�W$%k |
��x�ֹ�4daq�����{��/���U��\7������d���`V��~E7�7C�4	=tq���^��Dt����u���ˉ�ͽ��]�����	h���]�Q`�������}Z}�VK@ .�` 4?אZ���>�����t����!0��K���Tڟen����VN*�$�6`��|��"g���24�)vi�&4���ou3����!}��p�e�2%�;8dfK���5��� 9�h�2`���-�B.'�4i�<>��<x��
�E4��8@�݂ڙI�[��O�j�$+;@�l)���!	����؏�~GH<���$n���ϻU�?�/i����S^A�F'r�U3�X�q�؟k���ͳj�?����?�l5�	M���S����: {���H�g�Co �
�)�<B`��"aq��3�"�p�Ҧ�}�y;s����tu5�n�|������!��@����Y]�/N�6�д/J��Է��'�oC���5���.��{�r�j���Z LL�[��z�Fs��2���	
��unp#¶=#�z�uf-H.���t��L��_o�ɔO�A����Ȱ���R��B�C�i�[�}ƍ}_\�55f.�>�i��^�M���������U�cPG׿�A�4ǭìv��-�6���� <�\��N5�~��:��2��o�H��1)@�����7��9�i�XGY*le���g�C����[ܧ�B�6`��N:��i+��	��ko���&oѾ{T�Nʇ���^@�B������Dt�O��R�xu-�[k�d��&SL���#D����l�IO�P�C3�v�/B�E���4q�y����o,K��N�і�R7?"��1�3_��*%4��w����>f�t��/0�����$�C����D=��\M��2BN.�^�|�R1j��c�h�g�_1~(�M���4����?k�;��ϝ��a�aɇQ��fQ;S����y�y���PҼ���|bS�Ň+FwKv�,%P���0�Ӝ�y����Q��_X]Ҙ<m��u.�e�r}&����/(w7,k�Я�n<�lқ�Bz9=�t��N�dLX�,bg1���1�~p^�z��}~Y;�������m''W��g��������n��~��fN�H�&ñ<