XlxV64EB    1923     9b0���&QA��y9{F�Q-P�|ޤ�.���SMS���Z�4n�<%]9d���4b�ED���a}@��z�3����٣�W����QӭtNMQU��NUtU����oI�+)���1N0��_�:��W"��~-R�طx����je�z|odz��8�1��Q.ўV�*C���k+�2�����V(���E��J{c3\n�����_=��<}���B2��Q�dc8{L�$2pUW��|�B�zE�_<�:>dP8Q�i���z�~d����
C ��h{�i�ӽu6�E(_�,�N�*���J/5�KW�D:Mg�u��1���2t�=���:a'HN�$G�`)i���ɢ�wP��T�٧�Ծ_��cpu>|Gr�س�9�X=n�[H�(]Qzr����H>���#�Q(��<@�o����O԰��n1�Ԝ��6w/F�b��$���O3p)�RtO�߼��f������3�T��m�2寔8�Bw͍&~��fOM�!~a����0C��l�3�]ڄsW�0�O�I�M�L�B��qZF�\����;Q�:���8>8u�Z8e.A����C�j��ѫ"[�*�SC ���{ٮm�W�U��<c��8s�<O�~t����=���6��$��P_��1_��U����(�>�VB����Ԑ�-�4�a=���� �O���s�����f{���q�H
\>�v�	BW$�F<���t�J�yL�|)�I@�n���`�q0~�|�e�+�wpA�V�r���c7Ƌ7�9 )���ݮ�g��&�,L�v��������EVٲ��kp#�)(��C���+��%Q��}t��L���m��E
P�k��e4l?�Ś48,�N����S��<�(�c�U�����F���閧.�}�u�e�>�.��=�J{$��]N�#���G.б���.Yjj���6�g����ؑ��RHOͫ�Z�۾g���ۨ�90{�ȉ#~( �3�]�̋m��}�@�SH��ܧ�1.����(ņ0�?u���E� �΅��p�˰�+��kEvE8�쮑ϸvN�4�Z��s�Q�,�i��ׯ��F-fsI���4�_K�Cl�T��+���>�}��C׳>�I�����i�x�6;��_�!�� ��wJ��K߽Q�M�V@�G�4s��~ok<�銃���-f`����� /���vJOBvO�|GAL�]nb�*���鸅f�[:��w�On��q�ć�3ϵ�*��s��B-�1��r�0��!%3�ю���W��a�vǏx>:-T0�g�L)w�Y�3n�"��/��o�������v�-�w����4Zc��NOE]D�S�(�I�in�6�q>��Բ��L�Z��Q���������)�� ��ֆ���~��,,<�����OM��397n��j���@/?�D��kI먃�ī$B���6܋��0�v�'3�KX�t�&�9��6��c����+O�QiI�.'���(��Cn�$��	�,���~ 5��C��-Qa�݌;���Ζ��{�E�]?��/�]�#�=�<�$\�5+u/��P7Nd����D++tղS�ý$Zz8���B4��Vv�_��/�S?�| ��&!ŦIz.h"�rǘ�&ə�0y�`b��<�K�����q?�Ǔ�[�o���wO��{>���(yi��s�D�^oƇ��AFR�{���8�'ݾ�z!d��ψW�F�\�������gO�U
-���!�}0P�������#r�딉y��ʹ����qd�mw�lJ��Rhb��W_7j=��x�?�3n�O�=����*��]0��;��QPt�*�䟿K��̷�Lȏvr'F�+ҙ�wV��Pٳ`��4�ϑ	��K��UX�ξ�T_����j�0M���i���z22�W����<1�k��*�A�#����\�$x̖�.E��~*d���Y=�#{\k{�iڧJc�KP̴"�_�6ؤ�I!�*M$��19��=��,��s��e�,�������.���V���8��\*�YiW��d�,%݊Pv1��i�*+d��X-,~[s5\��~�E'K������X��?�O6{�_m�[l8mHsh��΄�{�v�����c�KOPK�Bū��ղۮ�m;S�?YN�)`� �����~�\�������D�V��^��t1�������\��脏��kק�~�J0^ܦ/�VFm0!�`�� ��/�<�:A���e��~׷D��<DI=da��ɼ�����*�q7 V��˜�&���.ݵ���!l�;���!X�7F#�s9������nHhz�;��!x�4��d�Y��X��n�T/��S
����G���ڟ&�!q�C�A��0p����!�P	f����kn*���c�������b�ZGTĔ�xw�̇vbS>g�