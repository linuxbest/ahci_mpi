XlxV64EB    1722     870����sԎ��.�o����B��`�������(K��Hg��ݜ+��D���$Wz��s�\w�����U2����b�0��Ǳ|�����ɧ�x����tXX]xgl�I+ͬ��V���c� �l����@g��T�[*�#I�I�ib�������z��)������r���M�(�ˢ/8�����ht`�7��Z,ᱰ�L;
�L�7�j;��q�csb�,1��)� �,�dG��Ey�d��{*$����H,h3���ҙTS��TQ�;�h�/\yXU}I��c#��m���|� C��syID'�-��Q��Rm8o���p�r*��GI�'�5Sv��g[K,�X����Dbx��`���Z �0Ƀ����RӃ\X�+�h�sbF�@h>�K=?£������L�H���|�ro�MhJ�N�so#(���;���)$;�!�M�M�o�@���q �̽~98�7��@gV�"��r�A��HX�Nx���6[q�-�?��YA4
�<�IR�n#b%�2#ew��#tD���N?Ѫ���WJQ6���	�S|���w�v�H|(b�ʵc��d8�CG�{�KH�C�JǢ1b���3�Z�����|�n�e�x����������	���� y�J���CVA�.�rFy�q�R>����=��aa����"+�����?�b��%���i�;Jx8��V��o$3��U֙$�׫O��|�i 33h����*a���\�f�Ӿ�=��c<d	_��J��f|?�S���[K�}b���P�T�n3-��J�)�HT*\�r�D:^��2��W�C����aB���E��q���!�Ĉ���ܞ&_$���2�t�#�4r�,��寎��#_SH��R��D���P�����9f
�6'#^oB!	�w�;��c,>E?�0�a�� ,����/����+�sh�f��b�o��P�OZ���VE2�y�t-��F���b��e���Ts�(Y�O��?$S����:��xej�?6���bqEr�G"�G!������Vz�Ĕ��'�K4�Z���7�3`��A8y�����B��b�8<�-���=�����<"����;~��M���<���ۋ�#��M��qxt�Ռ���<�4�S�.�<m
?��.�Y��V�X�X�Q$�x/z_� ܼ3v�:����8�Hr� �E���P�����0�s�!�����l��/"\vTc:�찺��X��HSM�=�vͲ�s�tC|��"DP�J�f�4ERL�\��t���4� %��M�Q��}�2�h�W	�ϡ-d�&9��k�3Z�rD�5i�cW�o��cQ�ȼ�g�A�h��
��Ǥz#�n3?ٚ�F���՝/�.�5	���m�3�[q�ͳ���Ư���H����$a��P%�G�ߤ>�*����yq�3��[{�I���
��i],�wG�m��5���fRGO;�P���Ԉ|�;͒�È��gRZ�e��'����E�`�%�*�L�;�X"�L�&Dk���4�a��ůGC�f|�_�JV�yz$�34�c��Cn�/��B�W���eDp�=��[�X[$ne���DA�g���	�e(Cy΋��r��ͲΘ�e��\���
XXcB �׶(�¤s��2��i5��My�e��A��,,�V��<�&RzB��EG��%��΍�^9��m�Z��z����󻰲�>�@ ��Z��Щ����N�kI�	<�WR�������KE7��'����3�`��~�L�GWs��+[_����������O���[�}��nŔ�.�2�}^��0��
�EM:��tܹP#��)ɾ��y��h4�z:�XQ�N�(��o��W�6���E�q�[���:��Ŏo2<�?Y~�S@�s[]�*�p�DT�!h�OI�,9M�l�čU�P�^��l�|(�5`�H@�٩ފn�0b�r�/��"Q�i�ʒ�
��	�E�F" Rȏ~�D��r���I�!9iq&y��O���TWX#�ʕS�9{�S�1|{�T���\�Maȼ��B��ֿ���]�M|�����d��f9^aU�����//�;�xC�^qH�D�'��/-�qa���?�a�$I�[S�9��(�KM