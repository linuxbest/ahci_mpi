XlxV64EB    25de     ab0���,Fw����aCÑ�(�[����VZ*7H��U�u�D���wةR�=;�m;�_rH��,=8C�k{��V"F��#[��C�}Z��X`{���e"�by;X�9�T0�6���R� gau�Wo¸+�@t5���2�]a�>�+�����L���yo�Ũ����?p�=w_����<�)4</��گv0�
�
t#e�k�L4��˄�݊�BP1 �2���{;6~�~b�����<挑6��~�%}�[x������v�М� h.S������@H�H�m�nu .`zq1/S�Trkԇ,0GD'�Q���T[xc��j�e�T�rpƯ�W*5�rh/^�,(+nu���Ko���SK�|�l!dq0	n�>��j���)8:*fM�l�I&����ɽU��W?d2�@<�5!YSjP �cn<�YU ��#=!Zk]"7���rE��3/�re�p$���Q�H�0z&D��Դ�xe���5�o����\�V;�ZW��A����e-�.�o?�V劦����}�#S��!>�����}�#ۅ`U�G���	�"N�.3*��%P*o'E/M��g�ih���I�q�U��Z߷��i>���73N��rM�Ȱ�t��0�����`;�~(������;ʢ���s�����?@+M���	|^�����CUmܛ��+E?�@�Z��	X�:7,j*�\A��J�(2o6b�W� }�^���-8��([�D��~lRtb}c})zD�3�ޕ������.�JZ/�@��U�r�Z�22BF�ѝ��9T��w�E 꺆�6k a��$�).��|6�@���WĪ̀a��׉��t�����%�Qc2�~�~��0�Y��1(yEc��������gCQ/��v�y����)��a�w�?�`/fH���NP�Y����k,�T���LGG�-���Q#��g.;;n�}�q!tN�@O���4�9x�rI�9���DMU�!� �`���uuT��#x3 �2���9�)�>�����&%@����-�0`R��MdL,�RKS�����P�)mk �Q<#��N��$&�3�p�	�߿�kM�������m�D�������;�P���|�1�A;��R��>�QS�(Mb������&xKIfp�n�.���w�	��Bϧ�t�W���^fJ���ϭ��8�BF[��ӣ-�9v�T�U-~�����MR��
@-���:wz�jgQ¡��6�o�[��[^��{;�#���?�z���v��0w��b���ܔBn�&��J�/#�I�H,����p���V4��������V��R���q���wu�`�1*��
.��T�5�� ×xvKg��!��]�k0N<��'�wt/XsrI}�{�w�ë�Hͫ��
�x�.�;ׅa��Um�z#\H޺	Y���u��2�(��3��UV��+*ܛ"Nbu�8=m�Ӊl��V���kD��T�7x�"{[(6Z�,��Y�n ���x���_�L7팡�.hkğ��ȸ�e���5�eߛ�Gަp��5Ъ}��M�	�\U׹����x��b�C~ucwb�-�-���|R����ѧu�EY+SP�06B4@U�u����i�<�ԣ������Y�?$�g83�{��n��X�_[;5f�p�����{f F�Xl�K��s0T�9��E� >��<�={?��W��㪆$�P-]bBT΀p��?E9��7��E���t��$#pw5�[8ɥβ��̥;�i�O�������C�Ab����6����<�Cv�W�.�P��{{޳�%*�@�{�F�$k_�D?�����#��eEW�(�y�@���z�g�S{f�p*Lw*]?�a�ȴ@�	�ǽ2�v�]^��ez����������H�n}�D�}hͫ>�{�(9ӛ?�]Tl��O��w�_�_�E�DֺCuI_8�	>�����j�%��U
���&��H�$�.�Q���3�o���@�.�;�s�)1���>Z�g�jJ��a��|���00nFc��*�N/��y �f�
�|�%x�Ä���r�m�rt[�OS5d
yW� Q@��&IE��I��78��ɻ��i�77>nI�>X�}���5W��c�k���
���)#p�p�u|���m�Y��+:������/�+�s\�U���*���&�~����y��J���,�c	��nxn61�,O�˲��rPQh����n�7�"8;�IQʒ>��X�$���1�;�G
�<l]?"������g��	-����;�t5�X�	kf�E�kb)��ɒ]�������p��?ҭ��AH?Do��r*c{kV&$t�r����sZ��N�b�К~��y���<pO1I�z�yH�V��ގԦg�<}�����%~�"���s�:t��g	+�� �^g�.�J���Y���0�>Y��ڑ;=� ��R)�x%g_�ԙ^��~�'5>k�r��Ez����f�I<یr�=�M�dՍQ����g�Z�kJY�A�M�d�<'�'΂V+�q��$u������ۓ�f��7�Sɕ[��k\&��e�~�X,�X���\�]D��C(k۬{Fu}'4r/��V�M����N� ��|R`]��?ooZ@�Ai
~ĭ��ۧ�)�"e��{�-�a���Q�} ��VEY)ʼ<>�P���L�G����V��n~m>�����.������ (ǫ�vʬ<i\�Y%r���[;�e�c'<c