XlxV64EB    3ef3     eb0`������;ti�/�ABӬӎs��j���#w�v���9���f7
G�a����Gaz���7�>����
՛�@휘��.#�)r��ꨐ4�f���p�T;'��K���.��G]�P���9Z���C�A�$��&۴J��%f�w�qj��?���B��t��	vW�ƍ�&�d�����Z^r�an_2�h��vBNmH;'W�c���O�2��ƴ�k�a��E���qX���F �k3^�x6y
�y+.����ͦ	��R�]&&B.�;hD316�����Ӛh���t���Z�+�[�Ϊd6��J`�"�WBe�NY�@	���&4#8�9l<W�+P��\��e ������6=�WyuZ�8.��n��TM%��,����q�(C���A"kS����9���#�rL�I����u�M�F���e��?
���ţ�k�Tݦ@`���g��`��#[Si�*=9|�����u�'J��W�D�5�6�әRl*L����(���0��e�;��c���[��G���Ò��z,.�O���1A�P�ˎ���؍X=2���D=���g��+C���Q��&W�?�麅'��ղ�dT�x8k��5������FZ��&�����,�Z|�^��E�=l{��5�-�M��;*����f��������v@Ǥ0+���H��L�"n�Ǻi�Zc���ۗ���$w�����ެ��;�۴P�idkP��g�v(�ˠqq�q��9V���D��F�'�v�B��+cY��O?`���̴�x|����M�$����L�����o@I�u4t�7����F�����M,]C��@P >�{�E�$�r���(���R�]=٠K��ׇ�܁�v~`��waQa$e86J��x�*a����ݴ>9A3'����a����I��l�k���>�H��n�N������%sSߘ�����XTOp`Wi��yI�D�=��ϳ����+FzS>m��&�	��d;Y��a�@h���O�� |�����c���sf��'G(/%����QR
�_�Uv*7,~���5��O�¯3�Ȯ�^4�Vl��J�J�H�}��-r����Y��7E�b�q���]0=�6Ln&}0#�Y�&���'�7�d;�"J�t�A���f����Y{"���ɕz�.bbr�h�j�:���Bkv�I4�>�����iBӠ��0;��NQkoٱ��;7��m���N�A5%��Nw�D�7�l�+� ����pU%U��M�̄9���?��-���j��y=���(�w�sܨ<����3��[��O����7�M�h[*���w�4�ccE�|Z��k��t"	ֱ���<:�o���ӧﱄ�E2��&8����:�
q��~���cu�pK18m���\�0�����T>��1lqշ'���â��u4DJ D�*Ƕ�M��*�`�Qwbϓ	!+R��E`[��]l#�Z�� �z�S��{��K 픃�f����z���`��ZcM��[�h%�^����;ox�J⨕��ܤ�P;�s��<s�@乹�M�;p����E�8�;�X4��9 g��@w�1<Gf�[ꩉk%�y���v���<HfS䖮��q1�>�V�}�'a3y��e�M�M���@Ft�������vn%y;~�m�!m��c:I�x5V�рv����v\�!S^��m&��lb�cb�,Q�<7����MŘ�z�9���`ӴY)ܓ~:A���շ7�X>�J�C��Mp8JzD�y�}b�a�Rt����?����j����T�±�'�� ���[A8�o:s����,�#{�bk��)�û��N�P�V��s���$�.W�1�c(�g�.�\,#��5Mik��9�,t-?T器�7o��TM��q�NnL�}��h�o7=�cz#N@+������/�o�g]>��Y����w"���>�?`������#4u�s=�\�=
	�mݗ��i�Ab��ӗwP��B��Ye���(�ZM*
�oW��§+W�cь���Ud�n�-٘+{�n_s��@n'T;��]�r�oS���t�����a���u����+E`�n K;[�f���Xf2:W�m��
��9��:Q����{6�y1�W�n���e�y�5`��#գ(����[� �D��^�r�����r�N�C��� �|��BZP��+V上���7��qO����V��.VJ���ͭ*�2j �4��:��S��9�6��p��{������_�|l�o�@)��y+_Ϣ@CN���C9�w���=���r�g�=�<i�Ú��[���
�7����b�)��xle�҅��P�m����0aH�u���Ӝ�<�y0ٛ����!Q�{�L�����'�
0#�b�P�Gxm�"<Z�_�B���6N�l#p�aVPx��k�-�ę��2���5oc���mޣS�f�u�U�I+�������/Ne]PEp\�+����G�F*xzN���U�X���gs<ސ����J�f���F�ڄ�Oie�^o���0�X2��f�;��usy�'� ¸WR��I�Ԓ�}�Y�� �̜�?�ڱ���x�37��(����J�w g��Ւ	�_vR�?Z x���}�C^x��zw>W��3(�(M�H6l�޿M�"�Joo?�h(0)#�Z��q�����'RS0|`�MW��W/�EެҞ�d������/�p�3�u��H��&.W��|[� ���c�&�-�ܶjzG���Ӄھ{rR"�_���QɄx-�MJN0� �$�4�Ns^P�;#��1Op4!9��O�,x��O^�)�E>5q$?������ ��tPQ�(l�
���{ݾe�Xz6<'���	Ƶj���a�5�d;�cf����I%�����xP��u3(n���F<��!m4�3�[� MW���T��_��B</���ލ�3�a�p�*Pp=,F�U�Q��ws�{N������<M*+����)-��2QG	�o\�xN�ѥ��5H�����U_���yADkݮ�9����m/���5xtXg�����+�1��Z��K1=���,���ʤ�����a<�U�|�!⧚� �cS�eTg!@rkU��I�c)JTqg��Y=�f�~��h4$n�a�I7"����حS���\o�t8��ҕą��?C9{�6�	8���Ϧ/���<���N�.�Y��H%�#��ù�~k6���Kog[�����.W���;�t����L-��S��0�&��D��-��'�z�����8��xX����)�$-1Xa3�_tC>�\]��՛E���*'�)+_�`^h����\1.o-���-��R��;��������fc+9��}���k����S�h'E��kF��N�8�8R6U�oKSM�?��~R�5�í��O �h�ے�g�`�oq��c���8{��]|��Ѱ�$\�Et��3 ���8ѡA0�>8�iTxu��É��)�<�����v9�aB(p\ec?�z��#����߃b���1]�R�]J�:�b�lIyAq���pĒ�8	�VX�~�
��tD�+t���
�*�Ey�)�^��b�K�Ü`T�ۋlS�<
�'z�%
Y�L�4K1�0d+G��%τ�8��Vʡ�kE�N�Y�$�h����^5��Q4�U�V{lHKA<k�l�-|�����ك�x�d��+���H�p�z@W;���