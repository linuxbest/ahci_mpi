XlxV64EB    1e3c     a80RA�H���jF�9�Ih�Y�.b�	����:_>W�B[_�M�#���=��q����!R;��3�ɥ];꫌Ju���^�����5����T�
/.b4�G(�])�\��e_-�荀3iO~����@Q�hU{=�/�of��uS��E~9媹%����c�&Y�����"���i?�g�A�R6F��?��@�QM��7x����S�ep��nk�CTa���J~����-�SL�}���� tǆ��IY�8����,��b��>*J��F�	�싇�|���������X�o���:�TW�p�����2�U)�{d��E�@�BCG�C��!Fg1~DV�Yl��#��M��<�
!c��8A4�f>O�	]�|��Nm@
��Z���En���a)�cQ��c�B��k���޵
�P�.iV������sGGP[	��F����Rv+�ۊWO�֮��z.�_������f�tt�Z�6p��[�V'_�|����=�f�?�a��i�]�c��"$\��8�0���gL����c`�e m����?^�.�5* ���@m��s�U�2�%b�����g ��ٟ�3�@.�c����	��&ݫˉ�Ln<#���ÓCϘ	�C�i�@�!�
YO��t`�Ԍ��$�5�q�p࠵��i�{�|rڛ�4YԒ��s^J��>��e�ؒg��ƒ��2c�p4{q4vRD# A�g`ўX|�Q�U�h	��3�ο`����t��e|_������{NV{ܘ��e�}�iHi���ZaQ)�X�r[u�J4hƱ��ʵ�_�I-�D�|�F~�n�����!mS7�������;5j�KJ���@���ЀS���n�-��()�]rSDK�7b|:���m��ꄏj�t�L���$��+남��FE-�h�bi����e<h���m��p��x��zVr5.�Ȣζ]a�3 ��~KP�jn��+SJn����g�s��"]u�q2��(���&���$�����L��8a8+�w�D�a`���0G�������QT�@�g�3Ӹs�U���R\ڧ��]�j�}Z��\���1�s-�Ǆ� �Q���~�w�:�P��M$X��5L�᎜��v�
Mf���,�<�Ox��-VH.��h�.��JV��TvO��J �83�k-�.!�K��w�,Jd��1]�t���*�����]ǅ��A�jJ�����^�"I�ȍ�f�O�2b7�����s�� �߾"o��}EVh�j��UM��pz��@R�l���o��nzkw.�(���l|����'M��OC"3��W.>ـ��Z�öX$�}(��`��A�>��ěʕ��9k���q�J��T1��#!EUK�������pe��A�R�ī����)�$�A��u!�/�u��:0U6���n���0}?,�NW��;�T܊[/;]�3���^�/[�b����td��} �^c�"d8F+l(����"��\ˣ�&-��o������/>f��t�L���c��T\,���ƭNv �fk6JU���h}�n�?.��r��0�:u�"��7
(�oх#�E��=Q>r!8>�Ol�oM�[���cNw5������E����ɗ���3�����>�� �։*�^�r+>�!����ad�jo���R�������W�A�*�`���Hu8RoJ-(Sy��k�wo)�-Gz�ȉ�4C���>v�_�<����� ߂�0_��������%�\	Q1�kC����k��&2}���w��ː�_� N.Jž�`���̬���\�9��q�;L&��k��`�2KW�5� 0�������2��l6�n����9g�S[O�Y���p.�nu�U&�zq7L��}�U]s`~�uj^$�d�+*s�֋)�C�������Yb�N��AwY�����?���R:83I�
w���՚��G����:(D��`o����b�y�Z�o���G�^�ӂ�|d��%���W���?N�G��a��1���
�S>54��D�H�B Z��b-��a�Owvl��J鲊�H�ᇕ耖^�@3�b�O~�^�ڇ��4�X`(Ǹ���IS��t�^V��fX!@�#�ir2�����d�9
D����ӽ��a,9��$�N�pD��_6�4�g�@�yW��W�n��1�5����Mu���$�_#nhQ��<�-��}\5�f1��N%�odG����8kEp|�"x�| �i�J�fΈ�J����%����NH'�������ot��\	V�f'u[~:Wd���ȄPp��RK��Y��U�P��>
���$�:pSԸ�D�DCf���	V�a��=�OmB��1�9�����p����A����Ƅ̠8��O���Oӿ
QWm�#̢�v���E��t��|��x)��;`G ��M�C���;1u6�%��n���w�� bWӟ�	b���(J %T4���71@�-�G��h�ݑ��>���#)�`Y[v�X;�\^��"ɗ���2�k0�#li�,+�e�*��X��x8Ȟ�,9WH���Ҿ�a��il"�jA`�.K�����^"=h���SC9�����G�n��)#�;%��_Ow�Vq�~tr�Z\���ʉ�,�Ğ��6�#��Uϗ��P�E�xM�#