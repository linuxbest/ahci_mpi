XlxV64EB    1fe6     ae0(���.�5y���B�n(��*L��=��I㯿��/{5&Ї��};��K�����2�8�����W�6ׂ���oڥU������-3J��8� d7k}�?�*�ܗ���l��68I\�r ���.�M�jI��ћj.!��@�Q����m�d�	��C���Y��@��HP1x@�_��s�z�!�}�U!Ak��{�Ds�`C�,:V�����;�c��eݷ�b��HK��:�P������_�������������u�g#5�cS���o�anV꽈
�	����\��>�p�%��u
������%x�ޛ/��_��7~k�pn�D9ar��-��WQP7�h���;r3ѐ
�8���"���Uכ���� R��!w�^�/cG��d� ���ˁL������Y($��w[�v?���ax�o����Ith�D�;UBL
a��l���XMqF��m�3������a;��i/_ܻR����E(m�K��^޿	˙�K"�z�r�D3
P9|a�O�4������Է��3��BW)�d�����0Q_R<�7'tyJ]gN��m�^2eH
��Sm���4&�@g�X���@�\}�?k�FX�3Z�"E�%z�m�)�|ԁ��zt�[�c��I�/M�S7�~��VNU�B��"�����&��\=�H@Fs�-��%g��õZ98��a���k�a"R"�N��P:�Ub�P������2Ny����@�m��mT��\�=LA�[����gƔpz�t]e_���t� f�\ֺ�W3T_��-<�zz���0�C��D[�E�;�����Jg�����-��ߏx5�x��M��s�d�����F-�  �(���E�	@�?�<6@�\�Eu�D����D�A�!����Z�"�J�� Ǣ�
�hm�����hE��*��v;�L�0�Vjd��`4�����Ztd��<���.%T{��řO��D׊���K�p���p��\Br喱>�V�'��6v2
���]�fTm�p�]6�!)��Ry��0t��؎�W0[��N&lc¬h�t��+��	�EA.9��̄*�1&�$�v��p9�5� �R�^���%mc	������#y�J�P6(��1�2V;��-�i]��TQ�q�~�o筯��C���������x�G� s��mfu�M���I��A���6�QzP��+x`���X �m���,���v�w�V�8�x�ki�`9��O=���	���*�;<x��*�{�uJiQ1&��Q	�P�
�A�f=6��jS��<g2/����O�F��*_k�k:�g��G�ܶ��YTt��Fi��i���K�bKL�oY̙�p8�6bۛ	��P3'CUB~N�h|�G���z���vX1RۜV��h�e(�Y'+��I��k��I0Dg���NT�'K�D'fa����y8h��^w�GD-ע�ھL��4A�ķ�T��d�Y&���v�~B���[�1�Ͻ��vW�r��W�e���U�lQ���M�!@�
��,мv}1�7����U������'".Л�!�v��DP�`oA|<��sK�B�(a�s)�5��]�0F���+;4.BG�li_⒞��vKi�� t�p��@l:Q2��-j����aI����+��Z���$��l�9,��#���IVh����?�=�ۭ�U����Iށ��3���פ�W]o��i�(Dx>2����rdE����q��2�yG�Z��T `BLi8����UWBs���&bG_�I^�6k � �	�9���=0Q�X��^v�:E���Ts;Mډ�Xå������js����GQ��:��c/�ך���˖$dđ�頇������������R��ٯ����}#-2.?��k��B��"����!�m��xI��o���O��7�����J�v.�H�������o�e��"~l�ď��f,R*qe����f���h��	}��T�<��ܦ3�r��;u�-��2Hyn�}�*�{;U�zO�H���W��� ���2KIr|�Mu�D�+��8���@�X���6G��{�:�r��	��P��������y� .�W�w�v��{X;WM2���H_��X�q �r\�}G^�� �4ƃxT҂��H���A;�4���MhMI�:V��P@��R�jCo���p9Pt��t��+G�D�o?6�=�B"jBW��>��]=��17,��|ův�?dஞ������R�87)k������`3��H���e��d��<Ռ%[�h�[NP�)�aM�Q���.��)�%
�&?�����-j����y��ܪ$�b�V�mlϸ��X9v�t ��5�^h����~�.f���5t��x��T�ooP�k�c�-����7�겕"?4�%������3��~���g�J������1c#<��!
��;��g��������4 (� v�(,�WF��ym�h��x�T���A#ąߥ`����}iq��%b��T��."6�����ޙ���j�`�n����sS��,c�=�W䜐@Q�ۦ�*ZY�a��>>�Axr����Zx*[eB3�Qyj���&�Z�+�]7u
�=�L�̵Ƨ��'��R�Ƭ��O�2Иk��#�\�Q�|9�d�j�3 7�rd�c��?&��	�DH¾��C�Xb�R���%\�̶,eJ�<��S4f�*�Yӌ��Hi�Q�� ��i�l�Ĉ�sFw�4@(e�	�AD�5˺�<�_����13�