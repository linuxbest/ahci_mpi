XlxV64EB    154f     7f0doe�� �ȓ&��{�@�g��x\.�����пT?�&�k�͕ec�4�����Wy��O�>��	�И|+*��R����P�6zS�H��ICK9�ؚz}��JڠF���e��R"FJ������-,1���TG��>X�	L��I
����~דw��d���S��7є�f���n�}n
B�����n���'`4zk�_N�B͋��o����ip�tL�V�j���	�Eq0�B��ot��_G��#o���atW��U����1�W	���.�%�b������J�-��c��#���U�eg��x,9���]CU�_�1�C�x�k����(�#�_�_�1�e+}4�%Zt��)�-�{��� ���7̂!Zd1+����W��f0��[vz
s�2tfB6��nQ��#P#�t��Zp�O=�����}�p��$M@�����q}�"���PCy��_*y����NI�k�(tO�lE��XJ���`;��z�S�ߩ��\�?{�يT�_�4i�d��NVX)��d�6� K]7:h&�[�l#�	��1����mh��혰��"��_Ќo��Y�7���<7����L�=�q٫g�*�|�sr�6v�M���ڕ[�	���4dCZ{z���U+�V�8�6��ǿ=4���y�[Ze J3���Q-�^AVy�J�w����D&���G�p�0����,��D���D�7���gk�D�I��޵K�G�Y����%�ZŨH7a�]u��p��zk��>N��(4A�m�P�$�X3WW�+��������ߣ�	A�c$U:����*Fe���&���fV���9��K��/8qUv���q���ꄜ� i���Nm�/`��F\D4�a�c'���s�C�`G5]e��{����42r�d�)Y�邼&��^��F7u2�ȹ|< u����ګ�m"�	y}�A�T.�
wJ9;־�y���e#&��b:��W����ߍ1"�m���ؓiЭ�:e�
.�%�Uu"�ϛ����n=���Y����~�|?¤4���#���WwIڔ�k?pP��aݚ��X�VR?�
x�����2l��t�\B�������$�CS�1e�@�<L����r��I��zm̃��(9(0�HS����-��2v��`6�:{�q�mZa��	�R�GFCmd��.�z���I�%��p/�� ���n=�	��u=dqtHF�r��a"|����Ա�{�`��Ѓlzx%�5t��l)xj��<��q�ꅺ�u�Y����b��RAA�t�J�W����uyW'(���#=V��S���4Î��7{7B��/Z�Z_��+�FB� �t���ˢ�1�Ou.�/O�,I ���R$dbX2]�C�������4��g)�;Tb;q��i}܂ȼ*/��%�Nl���L�U-�p��(�/����OV���9̩!R/�T�/2��װ���H�Q��M��l�0@�O�w�+�H "����C��6s[�mw����fup�!�9W.:gځ�p:<�W���-�m$�ˉ����O*���β8�4�� �E�t����_�])K'�Ӭ?�@}�^M� ��&*���[=�EU�N���O}����*��8�[h�
ƌ1r'G���A��/w�������PlU��Q�4�%���lس�@�,��c&�OL�'����kl�0D���B�r6'q�R�O�9��>��M��l:%<���<����5]ګ�wF���O���$D	ꟴp2uv�����������l��`�y�4���4�� y;�M��G��_�=��jU���r�pB1�@%�k:�y��D���4���YQ��ɐǉ�S�O��ƥ]_UoS6�y�����4���T��:��hԩ�����T��B'�7�o��s��>�f����&��|�'NM�A$��GS��� T*�>�XDP��CD �M[�M���]�R��O��B�sϺ��2��a�]�lP�%��WY��� |"R}o�;L���������'�֥��O$��B