XlxV64EB    54c7     ff0[�
����
�0���8�Z )��\H�a�/p3-H��>�J�����K=P>�;}gy24���TI�	��&�c	�>�2J�an:�f9��g�	���e�K�؊�Q������q4�d�W����*)�ɵ�tJ�y�Gx�,li���#7o���"�LF�:�Mx��\��.��dķi��#���G��"�������2����b�GZ�kU ������K�����ҳ}�����B�xn=*��8�31��*���.��+�gɖ���n�V	Z�N-1S��<�k�<ԉ����N{���H� ��!vómQ�圹�twZ�(�LϿ[k@ĝ����|M����d���dfEF�Ν�l�c�� ���Y�ϗg��=/��f�Y�>oT$g*^���F��O��&��9�A����qg����m2Ɨ��N8Y���T���t��¹}H�Y�oy���0�e[]3�[K�n������&�I�;-Wa�,i�{XQ�Z��^�1�0!K���h���$����Rx����{�}*�+��pEW|�K��8�Βx獉D��8��zγo9��u�w��v�O��|����m��[�=zG���F+�ToM~ږ��Ln!�'��)�ǁp�� 0R��@��S�*d2^�����(���W�Dn��������S(n���j����̎[-\���L�wi����6i&ڊèߋ)u��>��J�$�8��q=�*7�̰�nq�I-���*�x�1O
=����w�p���IBB$ϑH�ag�F����/dA�Q�������kʚ>w싮�zg�bݓ��F��%I�z&�l���F�Lm�0~8�6Q�,վ� u��޷V�n��Eј�։jF�^��օ�P�V��I��
\��Q-�������D��J��W�Ð�co�	i	�C�譬�p�-�;��x�Y�>���0Ҙt]H3���h�y?_D������u۹��bB K^2Y����|�e������ �"�Rʯ��۱*�1��2۵�<��+F+�7m8��jg�rȑ����e1����چ
]\EL;����F�"�%�_P'���v�����a�|���ێsՉ��������uW��pZ��.�%���q�W{�L�S�x�ddQ�q�;�p��8�Q������bF3i:l:g�h�i�)�Q�^���{ ��	�G�)|���a��S�Z��� �v�v���)�(&�������v������e��s�~(N�/��w=��������m�L���:��ݥ�X!d(|j�0a��/d��EC�}�1b�;��\-@�ZD��Lw�lY(d!:=�纣�}����u�����|V�D���u�O�#����G�1�I
��ˡ=�k���O�"'��/�08H��@�[�j�#�K�?���Z���+��EY�B3r�Oi,;6��A<*:�-��ɉ�[Mީf	��z���o�L��RC�h��F�q�����y[5L=GW��.đ�fc��">��D��A[�����{#c��l�Z�V��>H����J!����@	�F��ݳ'��o�󱉓�v�$ѿ�Jd��z��q�Gˋ����Q���\z�Zq��:.6;P�&��Gz}F�ș���M�+l,�Px�HU��
�2;	>�A\�� )/'m�C`V=�f�&�U��$�Ŗ�`2�9�����*2H�I)�!��pzp��o�bg~��J�S��z�KʨI�TI4�3"��� e����ʗۚ!߱����
¥�lߥ�Cl�'y���IK����8�N�Fg�,����5���a�o,M-���[�в���)�z��v�Z�ⱗ}�[A����9��0{d�՟���Q���mf��o�JS�i6 �]��  �ev�X�� ǔ��JiA���n&�o����P�f@ɤoHퟂ}T�,���,�,����SI>��8�T��?$ʃ��0q�¹	�1P+�d�=&�P7�&E����e��4tװC.cڜ)im
T;T��g�.
0Ǹ�#Ѐ�Q�9V������e��H�����Ƥ��%�QLdn�k��(N7�'�'U���k�RcK�oq�z�|=��s�+
�J @~KL� ����iPU�"pO���dg��O�P�Yf��H�!�(-�Fv��O�b��6� ��j���|b5y�^�X���\�6���0�?���MaJ\�?�U%��V�&�_9@��B|?�+&	"���ْ,b��.Dm��+����0W���ms�e����Zn5G���MT�d���9R׭��Ż�k�d&$d�=u5��:*�y��j��~KQ�#���z�,�]��b�zd��$i�����8�>��s���[����Y6J�%�@د�>7���w!�AH��7����ǿ;��2oɲ)�F�Ep�g�@+��J���?���'JL�W���B�>��My/���U�8E��֣/w�8�~J�{�s2:�dZ�[Si��E0����[�ě�}==Ę�ؘ��!Ց�����iM�ƊQ�u���DGS,���5�����Y���:�Q��Q���y0��:�x%o
��~�� �����[6�T�Έ{�)aN�f���;����,�(�����o���V���Qe�aCJ����f�YZ���IV&��]"�m��J
=���Ѹ��|mʦ�Z�8a�?iH�*���2��	3I�ؗ�!��c��tjf�`��X{�*b�Uv�||T< -]���@�p���lG]B��å6�2_���l����iY�N}Y��ԓ��9[����Ge�㋏�-3��\pO���@5g}Ð��5zt�MGV��a�1;�@9|�R�)?�K���P�|�^�9t������ݨ>ɥ����$ �f>��=b�7�W
��[�*����>���qK%�o��,����~+��輙��ϵ�$1��V[��wB�`�7M��H�(x�Cݾ.OpIq%��WS �
�I	�3<��5��)}E�Z�/��U���IV1��0�!�@BL����4*ɻA�Z��@�g7��.5$,5>�����FR	���Gj�Q�D��\+����3��^>Z�=}5փ~����V�:�����D1ǩn9�}>�K�:�L�w .3
Ӵ ����|ʌ�j!��8���ձ7��*?�襡�J��]9��]ǹ�,�~��
`�[���P����8Ӧ?x����;��B�%�=Ϥ_�r�:���wzC���ԎlpC=���s6g�q=�(`���&8��śB��<Ӆ����)����Uhr���"\p+����Cބ��9��J��N��#����M>��H�zX���Z@�!�ɻ��!O�p�a�1ѷ�	�k�gںX�Hw'[JE����c{s'�'ŇrQ�!(�,�0�?��	��
k��a�wθ>�м�t�(��4n�(r��E ��c��f�M)6��V�u�!����Y뻛vw�D2�]:|����8y�ɡ`�����g�*vÃq"���$�q
����8r�weu�/2�"ӥqj��>�>,����&E-3�B��|�l��P#��h��dpt���b4�R@>W�>�.�Lo`�́'#B��2�ݛ���,��d[�ar&��z��M���g&��u���<S?<[����am�i�NƗ�	ݷ��r�:�vR�O

C�D��<��%O� �}s�����8pB����P��O��P�~�y��j��W\���j���Ґ�"�t�BD�z�O謶	ħ��G�E��PVO�S^G~���UC� /�_:n���]�5�.Srl�KS=�����^�Z+�h��y$��v"M�mC���K{�QՆ���4��4�	��R&�{^ �v�Xᑾ#ɗ�����V�y�
>f��]N�_����͔�؊��@S9꩛#����R�q�Sy������wu�[��g1~�qX����c��B���7a�����4��vJ�]��.�O;#�)���K�=!3rE��8,�,����Ɩ"��(R�zڊ�5��dס��ϩ1�᤾�w��$�Y�U/�Ǿ~����AU?<~&ֽM�/�