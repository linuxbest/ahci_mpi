XlxV64EB    2960     c00���4�A�� � �j�itK�o���?o���lb�w���u�Õ8���X�S��vQ?�����"�	gb�����TQ�]�%r�/���3V�^�a�V�>�dU���1Š��PSly,�튏�Q\q�l�7�8�nwR<ϝ�
T	�a/WH緮�˩߼]��]�]�Q��hr���H(�Ӣڰ�W5d�"_w���	U</"(�%��N3H��5�"��I�pW�ă�A�-����̰��͕`�W�;���&��>����5��#D�τ��G�)�{	�rah<��]�.�*�7�P ��wGOEUG�"B���!5������Y��M�2]��m�����̿��D�&^���J̙࣡o�d�C$1���)�lk�����5��r��_?w��sM���)��O})��R��zHHl%W��[y$�C���P �G��@!��vpպ��p���b/[VA��Y����]W�q񔢥��&�(�¯�ᰏ�����{�N��U�,{Q�7{�CMp�E�G�Ĵ�X&ئ�#�<(ؘp9��}�9�@�-����Pl���a'-Ȍ�V�U�*�:m�i�C�Ĝ��Ҭ�~� ����v�ʟ�FtzWS���w���]��:��s3�elf
�V���7H��M���fjIr�'��y⏀�WX��"5Y�"a�Kp�_� <8�RUۃ���G���X�r��[P١>'����!c�e.���H���h	>�IP;�,�R�t����uJ�ݡ�c�)�$�r=%>!��L�s��0���#��',��Fn��I�e�j�%�1�Q� �N��S�v���řOe�&�:LU����
r�-T�i�N|H���/d�b)ژ�6��{bI�����5�t�)]�tm�ȶ��=�v��ć���pN���k�:�����v��lg�iϕ�GPp��{��I%�-�{S�[�e��2��~�Kv'���(���<�aj3R<6X�.�B)���/��p�H�c-1�; [���tUB0fY��[�QS�����������E��Ԝ��)y7@3}�ѹ)_
H���� 8|�����'��?)=Q����ߘ@K|�a���	G�8x�I��>��q�L�Ņ�b�3K6�E%J��H�I�)�N��-���Ǐ�ֳ:sD"u��A����O���r��~�g�����0�r]�/0D kd��h5;�g�`�w�
��
��!q����C������5��@��V'r3�y���4Z0;^"K_�mH|t���ך��u���-Ih��5�Qwd���֡s_J���ʴ\u�sP���W[�|��N����V�d��寔p;@CY"�$�Q���'w�p���8d���5�.�����2���*�9�{�� IAJ��o�6͊}KKG��c!�`KFDz�!��0��IO�⬷�,���(y�q�K(mѕ���j�t|���i���̺�4������CӒ+�DH%K��#��+F�U�ю߰�Β^�"��e(��lhX2Ek���As9qB���Y'F��_[0��?�����Qړ+ټ�0�O������s]l���K��6x�޾���Ņ��jj<�A�=]�Z������%��76g@�Y�Zxg�JQia�tʡ�7�n�{ئ�Zi4�]n�玳r��[ݕ��uU>�z�7�S��忳<e]?=���C���7r
b�^>/���8��!��6��dZH4���%S�
 �a?}�F@/�� ������	���۰ů�%d��PG���U��R������ϙ��1�4z��w�=&:4�!�J࿝O1Ώ�Fm���F�V�&��ɕ/Oˡ���	2��7h�Z�[�����=:4�>{¬0t\9#��iy�+����&{�c;�_7`@o�q�D/�g����zd[����{���t^�e�g�r�	�,���OW���a��>��Sp�S���ƹ�z���w����K�n����&�㷜0u${l�:L&��v�6Ȁ��T�D~����a�/�/Ֆ�v��
 �݈B%�V�%R���yM(J���u���g_1���<�,a�C ݨ�.J�R�U�-�\�~@�3ᘆ��T��BH>�6�c��O�����':*��y�����*� u�X�4�T�I�Bx�0�F�5]r�v�n�Z�]b�zS�mq˚˯ٜ�d`d�@9�vH�p�mFťZ5#1s5+��C8 #���5�fĦ�K!�o�P�D��\f����/����.5����+m\�'�\�w�����vFN�ot!h�忋�V�A��c�j�������!'�^��d��f�Lr�Tf�/0�X����`_�T����/X�K�Z��N[�ge�4�b^�����k$�;\Onkݦ��?����C)�Y[a��^Q� �j�wX�D�����v:kN�)�^KvGN�'���1W����ӎ�,e�Ӈ�Dl�Fީb�K�տ��0е�VS۶���wU*�X΀ܟՊ^�t;�/Ќ�4Y. J$=?Y�ITz6'�+|~�i�Rf��t#(M�.W�*�Ƙ��1MS��a�����#Gr�d��u��D|�8�/�^�O�[�:�.����EG�C��*����Q�;�)yGdir�i'X�mH�mZ�b��^UR=�PcY�1����\��2��.�޶гv���iP�(G�#�e�2С���r�'�jqe��n H�W^Jf��8�R������_]M"�.��mKX*8����\�e�j��ې^_ԕ���L�4�����s;�n:ŭއ���Cy��$����+�f��Χغ~�o����基���5�%C���r���5L���=�w���gb�V��C���BD�������Ñ&�k��渵җk�:�$+`��P�ᩈ�Ep�C+7n�&��;C){�OT�
^3�>i;6�=EKͮ�3��hb
�8���<��_G�uR]��E���5|�X�UAh�9�l�H�4H�;9#�~T� ٦�~k��ZV�L�E]�v9Z