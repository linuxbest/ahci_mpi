XlxV64EB    fa00    2b607������g�����ݏ|?�D�.�����:��S����@U�&����+��93l����k�2(u|�v>z�?��'~EmF&���:���>�ت8Q���AQ�q�u�p<��7�ı�͠��%èHp����HL�9s�&C°򬝮�W'�( ��;e�����{ �����Iڄ�:���[]��7��0�L��J�z�rY�&n�TH!�ԙ����ɍ��FLK����Fu��g�p��&��!���沢�����^�Q]�|��M���_����QO;���[��L%2�P�ߪA1WV�jrYM�N�l��3Aa/�����]���ð��jIsذ-R��K�`��2���(]��ĝ�΀���V�������������n�j�>N<�)B��X�ϩg;f��i�J��_xz��6=��3(�A�OL�l��2C�~a�TG����no�&���I���[�!U�
�;�����!�8��>��xr�jC?��-ݴ7P�i�\ZqR�r-}tm��)����*D����5If0�?�V|�:U�>�LO���=EJ�䍢�8�\�������37b��z��6��+-���2J$�S�Xa1��v�6�S�3g�Oㆃ�ec��^�g�n���h_y	c!��M<��[Nᎉw��$+�㣿 q=u�D�Km�E�&$:C�0�:a+��s�]]�Kz���I�ЩI��3�t6�C8��K��8~�]`��U��/Tӣ9K��˔�H��BŬjG7qv+��~rM���⍭�O�5P��p˹���a����h�룽�y�-���*�h5á�y���R@��  Z�w�;CSv˞��1�5�0����'�}�j��#��@8M�'� �[��7�4 �!.�*�.�{A�ɬ��|L����	�_2�a��a����z�����bQ�'�&�i&2�-n�yKT��c��ݰ^;�nO	jD�!�.�#N(jQ�.��`@P�t��9��ƒk����e�e��>�!B��J1�^�?Nmz���k2ƍ��\g�% �@�7�s��"��	m�߾�` Ӹ�Nk���^��d�Lj��)A�(6�l�i���=�����2(�@	�þ'PB`߁pG"��g^|��[�Vx��KN��eovEiȠ�\CK���J�n�ut�-yi
Z�)���*�׽u4��P��	���d16����/_�KI�"�u��� Z�	� �f��t�<,O��ޟ�#-V��q��|1�ʣ�_;Ǎ:CI����o)/h8-ޱ�����h��d������z�Bt��4��TnH�Uҋ�������q���\A���L��:{���F�)�4�j��z������.b&L�~���B���J��E�A] Ȑ�D�o�����<$U��R��mdl�ͭ����;������|i
]wTV,!�pz��xQ���E�W���%�N�W�/��|��0�w��k�LP��:x�����A+���d2+��2�)�+0

�TGI��ˢ�H�s�a�y}���$�pI�Փ�w�:![S+�Qޤ`J��%B�囓2�ՓH�[��8�G��|���{���i��T� O�~�'!?���بy�"@F�	f�0��¯�	��Xnq"M $/V�D/�٠�
�T��wЋ�����z�Wi�wr3� ޱ,��J�G����AU6�������qD��NSy�;Ġ�z�/P_�=�RTٞ�����0�e<#���(�t��q�����mYmEw�hp�F���ѫ��~��pm�ݥ�Y����\�����BwҰ#����� �=�w^�x��:~�M� �$]8��*Tn.�7Z.��Ԗ�i���씉#��pa��Թ�l�4[G�a�r�**SC�1z੾��U�gq�td�:����?3fe�?[V��;�����Le@�1t�ܜjP�(���-*����ԩi\2?�T_�}+)��_�]ĆM����6K([�fLhv�=��O}A
@�x��%��Ę�`hXr'D vJ�;�E.tl5]�2F�9r��z�=��o�`"~�`%٫~e93}ҝ�L�C���@rɶ|��d��d��Ѧ�fF(W�Df���s{#�`q�(nVAS����AS���������c��8p<�.ʺ�s��ʜ��2MnR���va�l����ǿ�x�� k<'<}��tv�aÃiw��u,���BtJ�mװCG|��y�T�FR-�<���۱P�ߓ�޼p�i�:��
������Ҋ:a)h@%bz��ʔ4����t��}��y�.bA%p��n���<w�'��d����مG0�R�]�K� SI_��,�E�2�蚚;m�p����h��(��RCVa]:�Z/ �28�B�9�Y�wu��?.���5q�%����>�/T}/Q�{|��/e��\y��U$��>?����҃䷭ߚ�ۖ���:Й�|�2�q��Ok���YHNp�!��G�'�b�����k�Î��<s^~ۤ>��3�B�m8�O#��qY&�P�j��K��mBzZ�l�F�O�+IG��w�huk��3�B��/�gJ�5kf��D���w{�>�gz4�}�5L)g?���΁A~��9�Ut/��2&���{.�>�Z_��$�:���>�G�͚��}G�*�,�3 �vfk���I�8�����p�Z���Vf�ݦNR9�M-�D[�"J�"бNY����$R�"@3��Pj�H��3BL]����~f"Wҫm~<�>�㻳���j8��ȗF� ���9��=����oǪ�R�(��|PV&�w�Ej�������	��M�a]ߥ�fl� "�I�:���_C����K�ive���A�t�5�f��������^��
G*F��W�Ă��F�z�����b�U�bͪ[H��0g���@U���V+�R��fY��َ;u��c8]�Q?��
'���"H��^�1�&+ټ�h���A��@Q�2Z_��<�z�MW)�~�>X���[�O/2�z����Ƚ���t�(G�[R�hhD@�c�e]X���H��P'�jQ	_vqϒoh*j�+��!����)y�j(p������l��b �T_��
�ۘo}'\�4����"·cT�
v9h�e�������~t7�\�V����7��0��!/׸89�2��V��]����D���C� k�|[��Xa��٬6>�+-"�d��ׇ���ͳ�Q*�.��"ɮ�^zCg�p�VV+��ե������d�Xu�SD/�'m��}�����<�B'���8�msIM���У_#+���j�	����&��|�'�R���&|��Նړ�Sk��v)H߸\�@ުT�����4�=t2^�٠��9'�PG#���T�q�b��P7'��y���{c��u�����@ ��>�0 �H�Wʭ������p7�jڱD0!�G�e}y��� '@N���r#�����=�s�Ο�u:�����z[�a.���=�	m|�m��>���
fȽ�(�S�'���L�s�t��+`(4$�{��i�H]�6q�<ۙ�q���V�?�d��x�m[P����1xF�0gH)�C�����S�%a����LA qS.��m�3�L��F\'�Zw���^�t�R����'[xJ�k�yW��ά
�V��@����s�Y�ƟT�Si-�m?ǎs :���f�Ţm-s��Fp6��5sN�����,�m�8a�_��;�$�X��w{Jlr�Sum9}���(����G�*�gDߩnݶ����H_����a�)���s���!�G��T�%�M/��I;���D�s����r�l�4����({W���sE ���<0h�M��8��^��=����0�m:jZl��I��4�.�z3H�BB ǉ��HL��$^�z��U���]��q`F�+�o6��v���dn�-Uy�ݝ)�����&�#4rS�?���-o��.���hΗ�Y3�N<��/����(�ѾW 	5�(%��~��O�67,Â��*ft7�<���t���@tYv�%�i��?���a_�TIy��i��a٤�Nѕf`;jB�=d��m�M�X�քh��5��?������ϗ,�~&��=�/`�\���
�x���a����5VnE}y),@3�K����VӔ�� ����o�a7�/�����s�0�y���ˋ�A)Z�8������c�I�A6^2'�U��y5�X\��[24a?;Eכ+n�9��&�u��w9���Bi��;&6H��X�{XV��ػsMY���K��;�N��T�(J�y����g�=�_��G E|�IX������]
p��Y1������V����)�����"��B�74H�Z���$	�Tu�d�u�U֎�S�W��v0N]K�&+>�E�tO�2�~caPQu"�+�t��:X{8�e5�t�F�'ٕ�Ɠ�Z������N���xb�Q&c��)~+'��tQxT�vٴ	�X�h:����`Ķ6.�@����'V]�$d7T�G��Gc��R��j5�,*�^?��QU�t5jm�����.ő*&����5�4u
[�T�R�@:i���[1t����5���d|�	KbD�9�:��A�65cs������E`&�3�;Sa'�ڶե1ˇ�t�0,Z��Hb��&��'��KG�5�чX�S��LI�� ���պ6c�	-�M�!�&�)�Y���+ξ7ϝW�Z\T�7���.n��)�i{ ��b���hjFKؚ�l�Lc^�1ј/5���.�2��̘�V�B<R4�"i���:/#^�.IZP�J ���J����!�Sz�\�.C#�$�x	�)�S�z7�c,��D�}X3�ґ*_��r�\e>&��!Ɇ��>k�H���n�S�fYH*���?Ǫ����8�m�k�Ɣ������"�|�����t���]�p_I�P���֣	�'up���pG3��k.?�p�=�'��NU�m���.�T�����b=XS��D٠>8��׺�Q:����1�w��AK;%���S���!�h��L
]�qK5���rF�;v76aI�����j�|\��0E�me��c�뙒о�*�o����<I���3���93m?ok��(�m���*@fǣ4/O�~�C;%ٺ롕T��2����P/C��؇]���BB���~�|_��8`5�#A�o�Dj=�U9��-/�pm��1��e50Tw���ʸ�g+[[�݃s40�Jܠ�&�������M=�w�Il�@$0��šj�8Q_��fd�?fX����-����#}�[Ԓ��T(`��T}K�m�S�3��O�{���*֨�5�3�J��cY�h�!�� ��)`¢�!��gdFv�H�4	�3�E�����#�f�r5T��MR��^ �����qC�����
�g�@��M�'�*M8�I� aCO%�:��M}���n�X4Bm��jxxA��V���,b	��K�Ce�gE�{��F𼡧	*X���)˖�K_g�:2d�#wO ��7���s����/W����z.T��?l�JOitg��Z^E���m`6�d��F/:H�y{٠[�IvF������Y�z�w!�+��m,��v�2�)[C���n���7BRI�Ҿ>9�OV1g|Jy��y����@��p�<����@����҉�9�زqt��VYS�	OgYT��ޣ��m��'5"����˶
��Q#�[�,a(��bcc����(�C�_���G��V��9�lS�$jnm5E��͘� ���Bi�����Dq�sL���c)^����󡧾�I���7��7.�{�Q��!Q�	2����-�;�}�w�V���h��-��<�wn���8������9+�Ej���3��2��TW;�jdB5��V�s��y���H����z��i���L�+�?����4*Q���u�^���u�~���f�5��徑e�ߨL�	����1bc�H�ΘĻP�&�tvt݃7�0���2�T{��=p�\Q��T��;	��噸��Nw��
���	�q��
�y'� �Xy��eb���E���kP�.\0KrKJ_�,}�RnH�#���X��a�=*�x�Iִ�DE����1�6s��g�L������XH�%���5oZ�6����l	�������Xy�9������~ScffNIV��}u�o�]�-K�@/��ih½�W%�g������#�#e�+r����O��ހu��͍|�'o�Jj#mI����� ��$���'/���x�����jn_3_>b��P^U����=b����݁�l��~3��G@�s�����~W�C��O�*�(���$��8G+�=�'?��g� "J�}�{��I��?Ӏ�-�m>?c\<����H����'��S:ڽE4�!I2͏��-ǔ-��F���S����_;�{�%���X�ܱ�ʇ�^c^ea,A?���:[(TZ�'3*���^ü-��������"	#�|�:A�gF�\x¤����$��a�O�.�DX!���;X<,U�|���{��%3�HR6�3z!���5��@�e�Қ�Kekj�3����&��diGa�-�po�����ܸ��b��BV̰*��Vs/9���UP��q7W#�6���to��v1΀�|�� 9 ^�->x%#�ס�.X/�����S��PüPq<���u^pN(�����n3��|���7�~�F��}xsm���5���e�����/ 1�n��y9�<%��ˑ{��/�#m39���R�BK_y ]6����a��h.fB��ڱ��炗�w�ԡ0va��)]k��c5T�	ŰϤ?)L.��������+iy񣡠��Ea�NC@%����6���SV�w�c���)��`GOZ6��6�$��M�ķ/�Ő�S�������.ٶW���=Z�Z�zn�T���M�KkCs��(?�>=��'��>� �x%���
�^I
�8�}J�,shl��j�E:\o�P	�,�HF)F.J���_	�oƃ���ٶ�m��/��������E�d>��jxP���K�ԥL�!�҃�j�#��R����Ɛ>"���P!j�֖��֣��͛!��~�,��kA���<�[N���k ��}0�dM$ru%����p�&��*�.�A� s�?�8���^����uE!`�Lkp�,�/0�E
ȡ4{���Q�"�8�R�oH�� ���&��+c�s�B����cŕ"��,�xC�1���Yɥ���I��
 x��!V��H��T*hJc�fm�&7���������x����;��cO�ma�^)������?�Q`�ą*Y���gM�~�E��5��]G��Č�]����HUqŜ�LH�wQ���H�,m�>E>'.A�b,D�Q��6S�U�iD"��5��뭄�$���W�?�Mu	yP-Ґ9��d���G��E�b��Hb��Mp9��P%�����68�.g�` ��6�=wv�����3/�7UiF�A���޵W�1��L�ܔ���SN.R'p L|h����Ҁ���J�:#w�/��Ԕ<����"}uo�cD�9<�^m��W������RDk%}��0E�6ϸEb�������ޞ�4a��2{_jF��8��*����oH*�3��AG �X�~�ܼ�7L-�%e�E�L�����{��,p1b����2Qf-N����C����K��
0l	O&��3۽�O���_BYe34�C�]��n��ҳ�ǚ�>	�܌�pe��xa�;��[�R1"*�ܵ�R!U?Ks��� ��|�y��<B�f���T��6$�j��C�d��k$R�����F韹G�'.�����ڣ�p�`�f��s�ٳ���C1��zP�|��h���
���}��Ι�/�"%�6�*��N�%t>Us�fX�Y)*m�?�d�nO|�-DI$:7�(����O�8�^/^i�Fx2�A��!&�m�S2r����������;�3 ��	�(G�T1�*����N=�!vƌ��ѣ��)�����������q�ߥG):Y��v�K��(�z����/'����=��4r��^f�V�o��4�Y�1��kb\�� ��x��N_Ǣ�L���i+�#>���������j�C�9�/��� �j�A�c��o�KΦP���/���Dp
,��ŝOH�j�p�����C��E6&8��m�m_�����ԘCi�wHZ6%�D�N���]�E� ���+�Qw���Z�+����2o��5X�h���
��ǣDye�--��,���E?���E�d��q�0��|�]-X���ʰR����i�W4�:�xg�2zς�� �p�-�;	�2���#?�B��^���˟�>G-!��#_/�w*EP�P,c�bm��{����*�P�D�	`eU&A_�0P=��$�q�+T�<u\wtz��xMqP��?�״ �̙��4-�(�;ܔ*����������A����F_��t��U������r4S�{(FM���S}�v�!��8�E? 6��GY[%���'T��#��q�G/���L���X�Sݕ�O=��_���\��%Z��I|nʦtn͠��ߗ�*�w�86��<��P���_��e��=�]��f��
�A{��2\��ڽ�!e�~Y&0t�����+���u�-E? oU��y�	��&w_²g	�ꧨ�Q��W���?�}GB �y�^޵���L=@Yw"�,^�H�:�w�È��B1U���u�[xV Τ�8�F�qK*���Q��A��s.&ȏ���ԓe1���]څ�CBu,n�N|niL>��]Tz;ut�h�EC� �|�����H��a�!��Lo&4bzPq���Q��0Y<��.,�7ȕ�X�>փ���*m�c7\� ���j�g�����v�;�g*I�3���$����y�z��z#��#:�F��ŢN�$�b]V�V�r�)��͸�m���
�1���}4Vގ� Ӟ�`��g/x���,��cK�&o=c�MDd@�G����_5f2�x�d��Ō�C}O78|o���(���b�s&.�$Y���G��+Í��ܟ����#�|Z�&ǂ����F!���>��0�����)�Q�e�׹i[�[�Ͽ��~U R>���{�ޘDl��ULm��%[�N�N�������[jeK��(�����s�W?�_�v_1d	j3�9/�S6y-�3�c���� ��es��ay���+p:���3�9S��fNvp!��Z�x�%s/R6�ǡ�і�����W<�xkq�g��@�!���kލ��Θ��.M���P�ʜ*}��ܯq�>0�̑����V��mBd#���*<�'{�\�7`;�P1��Í����L�<�X����R��4�����'��������1*R���'����C��0�X�qVK�8�$���*�_T��Z���y���lv(�-���e:^r�� ��Ĺ=��: L���f���ML�V�}V���8��R��J���Ě�����3���>M��!J���V�&��o%;5W�)��@����.���I-��"yo�.�мبЭ�-���eC|�~#��0N͖�����ԑ>m���(`�'��O}�5�<��I0�������l�� %}B�qCQq��:DJ�Q�C�����9�r���N�<Y��ޘfu0��>׍=�k�1���G���-]!�A�M
5<F����h����
Kia'�y7=�_n���w�X�A�i�[m�8HE	W��ۏ:݌�7'>
�lb��;�d���Z'��IF,]�>i�_�q=״/~�d�*��,4s���u�(�C�	Zd�"��@1I�Ӹ ?�=N������i����X�,�ҍ������Tk�Q�Z�pG�n�$��9-�9��x��s�x��$�v&ƧO��L�
b	Zt�i���:�Քa=���t,Q}�v����3�]�8Ʉeq.�׮��U�����I�� ��y9��9���#J�l�Ӎ�j��e�h���`�NE��َ��Z����#�7�R�l:�FKF�j��1A���E��!�6D����
5�)}�Ö=����4P0�S.G=6�c�Q�ژ��t;-�GR*,�B�*�"���ʈ��M��U���*C�q�}b	�)K�Z�	C+H�9X\�}mX|K�-R�����qqXW�GG�݅���QRi���̲�J֋�/���q]�1Y��@LJ�wR-���X�C?zȁ���4�L]�,�)<����<M �8)�:���$TE,�\�/��8��D�޷�w�ӑ<�o�(��s��__,V;�#3�j���R[�����+e���A@��W��%yN�M}i6�3��x��W��n��po������j	�B{����i�m��z���)�%�esgC��&[S��r���R6�Q�\0�z}��'�M��3�j�.�/��]�P%zn���E��U�f���$�;�,���埉ܙh��_7Y}p�q�Є��_��!�0w<�F�{�
�cnH�������obؼ�e�*$�h��ܻ��ɦ����z�ˤ	X�c�� �x�as�/\.]�����h��
��O�3_:$�J�A��rFT)B"dH͇�)�cf�'��E%le�J������vmxr��T�^�}��V�։��c��ih�s)�����J������c}.f����f��D�!)���l�i�p�W�%�֍U�o3�t�5��t��L�S��p�b�j����̀ȾyO4�V�F)�ʱ��g���9���P0�ƶ�C�T�	�� ����N8��X��S�l��6�*�.�ruB_X�B���#�޼[%m�E�#:�Cu�n&l�a�)��ڹ��������(����?1�r����`�$��m\W>��WI-N����!��{���j4A��䞎�*�n�@������p�یy��Ǌ�5��1K��� ��̏�j��j��j��jrXlxV64EB    fa00    2810�L!�pÓ3����O���꓂���tjҌ0Yvۄ�pfH̹�c���+���w�H�}4w��o87.:@}ԙXs<�EqP�R��/U-����͹���̻rU_I�Fy֕���j$��{`�妜A��--��ɹd�2��G����Y��V� ����u;�Gl�BIo���}Z ��T*H�$FW��z.�����**��M�?����{	qP�I�d�
�pܷXCϦ��^��U��$�\��U��p�؈�|��78�+,���jo>״�S&\gL8`�Nb6$����g����[�$�ce��n̆Fsѓ\�xJ�zH����ӝ�����y�8:����4��8��U.b¾�Ǌ/��|i�R&�RPT�9��#+=�h���r�vv�	7QD��Wy:��0�Cq-,�d
��5���'�)n��*C���+�5��ykS*��HLF�{!ŭ'�TW.�@��#��USȋ+ܜ�x:��8A3�au���W�)��[H�ut��N��EY������(N��gN��f߽/�;湳,��>���b�Ԑ�I�c�P�@�h��N�L�?��'� �����vir����RE���p� d�����eV������BM>�5�wn!0y;��O<ğ�^�̫3��bl�eD+�-oρ�Ǎ��X�e��|%��@�4��׎qim�)W�꾺�?���feL��N���>�N��]m�sm�kSB�s`?`�
�3 ��{u�i}Ѿ�o�뽋�Z:|���;�f%��j Q'�
�����[y�rr9J����2���AD�� ���BL�##8�dF��^Sb�:x��c�����v�ˆ�*i�rȯr.P=��� �i3���N^���،�<��iǅ6��r8��%���м�ݢ/=�X"�?-�*�PpF��w��LZ����T턲�B�"�S�w�^:9�F��Efx��w�m;	P���V%Ai'�_��?�+�����9�)fe,�NA�'.�[$9(�U����ѐ�c�C-��faB�"P��c��pN
q��o���Q�
�����w/I�LRܸʁ��0�����މA�Zg�l�|�a��#`����1�A�1�}!�-���|�{X#�X����!E$�7�ܰ}��i�Rk�Vl�2P�
!��*hmG�\z� �ԍ�<�0������1Xn]Vk�t�jy:ϓ���4�/�Иؓ���e]�.<�U�Zꮨ��;����5Q���4#�--q��*<h@c)�����m��gM�"^23�r\��M�#��Ym�C�q�RDY�װ����W�J�Ԛ/.��zc��f�X�s&�+�
w�:�
�m�� =�C�Y��l��`P۞b
=l���Y���E$��k:�(	WP[=�T�j'k�I�6��<Sk�u&��H����b�1>g����c%�]�a��52���C���v�vD1��)�	��,3���]���-��so�3:�އB��G�O\�a��ǽR�Zw�FF��ˊ`� "�ҏͦ���(��4;�X��R_��-��MG�ޒ?�����[7��76H�+�*݄�F��T�0{k
�lo�'���o�0��a!eQ=o�I��{�֢'�X7׽IN�@�D��8^�<���>̈#��Ig\l��|��&%g���k�,�Z����bފ�u�nn���J�^�dR�e@Շ�n��"���HZ�5�ܭ�5N��f�
�6;d�����Rf)V�ڲ�Q[�I{I���ۃ�gt 
��~[��<�bNHlI��o}-&6E񶊨4T���25�h⎹��%�y)���FC�"���Y<8w'̒�Y�$������0B�3�����@ҏɨͲ��zĘ$-PЌ�^�N��@do�����U�ʯ���n됖9@o8t�$�ޤ�M�+ �Iyo�q�'�%@<�G�n,~I�J��+a'��ћ��zH�U�=� ��U�^�&Wx��)��c�
Xs�.�K�W�_��
7����eu^,��@���Z
˃=^;#��z�5�.p7P�ޭ�<F���Jꃹ��{���$�E+�>�D*�v-3��=H�_�����������^��~��}p�̐H�ϴ�N����p$����/���_󄿛j�י��o[��%O!x�
�׭��Kz��������������!ICd���;��<�%�7��o��?�� ��?	����)�Q%
��W��Q\�|�f*�T�-&g)��.�����F��pKH�%,=?� �(�0@�X�e#R�M0��F��S嬹ժ���$DU�G׆�t,� ����͢d��K��
��<�j�5�S�7�PqU����F�){�zn��g��'}�#<4C#�����X�嫆�%yB�PP]jk�rj=���C�� +eݚhU:g�Nͅ�<*��R������(�	1��2c��p�҈�b�Q,��_u��Ο���9�We���-<����V�o&^m��{~�kcySe��_�9Vj���*�x�(2�&�� H��~��Q�`V�#�u#���l3BT���W4�Z�?Ea�_�E	g\�FZ�YZ�w�n`�����/�2�z��o���Қ�(�R�9}�^��]p�+s��=�M�uƷ�xo�*V��3���(k�� �K|���}W?��z�?�s���e@�"6����4)}�G�"�G ^B�, hç6�0E���|u�I�����!� t1h#�ϼ�_83�[�g�J^��H�Y8_��E�<���7�����7�F�$�S"�eE��@8���Xy-��N���F��=�+X$�snx�� ��~5}��ĵ�_���<��c�+m�J+��ϸM�ES}[߷��ӽO��	A��}��G������D1͓���RL'�*T�7��� ��H�
�����L��d�絜��8�w�C��ϸx���s�O�^��p��}��H���r)h0�YW���l(�#8EE�2>�_�oW.~�����K��X�а�^{�T,�8y�c�n����Z�?�LG���_��.�1�w��p'T�г�]�5��4��s��9�k���M �^��&-T��V���$�i��� �D�wc����~�%`6�Y���i�SR�a����J[��7�z��cad�.֤�CO�m���W��J��)�g���q�d�-�[�}]�ǩ���T��* Mk�򻪪�̰��\�z�3�R�zA�σ�]�nM��[p���j��.�%j6��_G�Tt�缡��܏�z�ˊ�Z�'�-��`^�C��D�m�ʄ��iU~E���-U(: V�C͈��=@�U�+��c\���onUm�	3{O�<�lGs�;>�Z�4��wz��7�jA���p��h(ߡ�O�ExJl~C�����sN�6��M�5�+�8�͔k�G�E��EF.<�YI���Ӕ��ps�z��G�|?}�Km�꟝8�r�	ҵ���-�_8����{9�J:,��wϛi�l�����;K��E�Rn�e$�;�e��rҜ��ʆO[>>C������Z���
ͧ�1g��u)��2�6b�Eaݕ���s2a! 4Oj�T
w��Z�}���'9/ߡ[��Pq��$�28�����@agz�qp'1�)ͨt��\nK�X���ڻ�R�Y
*�e6}m��}nlT[����õ��yӘj��Ǿ�*_'�w�k���OڔW�겨4�̪)���c�e�q�,�O�_`U1&B�C�;�$(�#e� E�g�,�UT���JG��6��k�A�qt�]��I`�;�3&���G.pU�Q�	c�ʗ/���b���#�g�#6:|��(�s ���ۏ�`X�|t�a�2�d���bٿJ��Χ��� L���64�����nJ�y��T-P(�Qi�a⒲��knS��Ӟ1ޔb��k�K��������\�k�h7��Q����/U����@��+o^�y%:VW1=�f��׈5	q:p�v��2vK�"�f�I<�- ��6;휇���b`N�}��0�@}�>��]�f�71<���#��IX��R�/���{h����; T;�9�U�0����'���ڭ]!�ǲ�C��W��"
��	�:�S��� ѹ�{���*�����P��/��̈Y�$�g<��Dc1�Xn��UE�})�J�_X]߉��$��B��ϔ��{�s�dO�-w6�#��患���2t���Q������Z[le0�{V��q5��E�G�rX5��׶
4mZ���޵�yH��h�fxՆ2���Q��	��\N�Eb�_k���\W4�xVvm�U��4��0�5E�v�@U4���)�b��Y&k3Ƿb�w�Y�z�C�D5����ܺ�iL�E����%�o�������|��fD��H��'G���L�L^<�V�������a�70{�`(X�
D��L��'_D.V���s
O�|�e^�"��^F<�|����Ut�;bKB�:��kɴ��tA��3�{���n�(^8�����%�{�'=�G6�,xCDT7O#��/̢�^����B�&%���v�\���=[�Lrq��U���A<y�P��ZB.�����B����/C|�mY�{��(�%2<,X���E*��rT�<d"�����&�4H�U��#:�w��0	�T��nM���@,��KO�qhK�7�PL�%��tʻL��һEL�Ʒ���5T*r�����2�ЅX���ġ#S;e�;t(��]VZ�(H^l�G�{�ﷀ�K���,q��C�{��|�|�FA4m��O���뼬�0(4r��t�rT���Q��Ab�������@�$;��T� W��"}����,37ߢ(aᠷ@*^��p=����x7��z���v�^���vPڤ y��c�BѹWH6Ы��`�CQ�+���fuM�N<@��8�R���		�rk
^�m��*U�s+u�׌Q:؎\S�hb�__f����i�JL�
�Af�X�y��C�q�ԟ��NLe
��A�+�t�[4��f
�,�������N��=�
���Β�\�'y5����a��8޽�S�\� aR���!E��6��<o�����,�a< ��?�:�����g���>#1D����D�o��������=�?�8����n�	†,	�����z�����)�v�1���CH<H�p��;����(�@�Զtd� �f+�\��k?��~֙ET�0-,�Ѫ�!�m���+r}�֫M!eϴr���}%�i����7���Z�{������=�=,-�� ������a�����U4�,%h>=�p֘��#���C�-Xڰ��8�h.��=6H%��:�\Ԓ௥��-��LQ����6CY@v�<>�  �L���ms����yH�uegFWW*����'{�:���a�A_�dx5]���'sw��8�zk�_�bg��c�*� ��0=c�L8I�H�/�0{qԑ.ip�I�إ�'�x�6���F,��P�꥗F��;��V���ۏi��_��$*�li=̩߃H
�TyB�q֟�4@
��2-�y@4^��q�p��A��؂��r{��G����P�2�T3��2��.��;Է�ߍ�%;'C�w�֭��XP�3���2�AAތ�[Ģ�a	�mEC�<_�O�j/��|^�:���Q}��Z���L
lF�?�G�v�����.k����?�g��CC �-��sc�߸~��8$}��X:��3���V���LM.���j"���-�4����1$�Oz�M`�a�C��1��؃h�&�@
��&Q��Q����"N�Nʥ��h���h�i��@wm�Ɩ�@�f���}�{���bߡ'�i�������������*7�3���C�b�N#�4�����ݨ
9r�!�s�Op+iS����~�2�r�ՏA (@,f;�,?v̒1�SJq�d����ݩ^l��Sn?�|g��9��nʺ���h.'σb��y<�wAY`51���=gqB�����x�-�y^[S[��Ԙi��M����Ge�C2���[\[��`�����U�aT(���\�l��P�j��j������T�z�	ѯ�p�	��\R���D/��[�"��x�V�X��z�y"���s�~0~�ԗd�W'�ȭm���������m���^r�n��i��ϸ�1 
6�'���$���؛"���F�)���B@�U����;�g��.^h�z-i]~3#G�L��?��w�\������?���S����:F�%�,������Cs�]a}L.�.�^�3�/ɿ����d�xb��屈�����؂А�ӌ� H_Ax��x�̊�j���3�|͔�S��Hv�H���|֥����r>s������g� �p�b`��qzJ��7j�-�����G�	G���)L�S�2��g	��!%ZNY.-��~�ٯ�jQ������SۨƝ|�_��{������a���;��X$Sq�va�0?���u���U�aVxN���8X��u�a�CU�=%;+��e[pD����B�$
���BV�[P3Lwu��zgj�M��%���r�!v�ǵ�,ݱ�G�-�r~N'���0,���&�K"�߮4�&�p����K�k���l�ׇo�PByQU"� ��&2��?4�{��<�:���@8�v�0h���B�"�+��H��Wx��Ҹ;���F�Lpm�S����j~�t�X޾�\��I����`�WhH���"s����Dg�U�;�����U[�}��@���>��&�Ei�m@'T!�%� �d��?�C����Rh��^�ɻ����#���ERօ]���a�g.te��G7@;�� 5�1�=,�=";�O9�^�3E�F�j�ۼ�L?{�b�)���~��˞J��GT"=H�J`���jL�E�kdO=�����)�LbJJ��GT2����QHuw�����%6�3§m0�tX��q:g����B8��*]rU��V��T�r�F�iW_��Y��n�����&�� ,�J���c7G����vϛ�S���|)�V�@/m��{��>^��/�c�&�#9�Y���W@�^k���X�
�$e�.R�F�
�o!�"��U�[�!]�I�����#��[���[=���������$"c�`omm�##�p"HpN;_�ÍMg,��^P��6���/�2�R���ɚ���)�O����8zf��G���[0���PP�e|NnY��(�@�h����@��_ϸ�$�^����գ����4G7;+r�R�7�rg�g�y���3�(�M��;L�I�W%�����2<�b��6%װ�����C�X*h��c%~h��<t .��˫������Oo���z�X� �>1�=���e�>8NW�+�lgf*�F9Ic#��-�)>Y~8��0" ˜M4&���Rױ},=L�]r�DN��K�A�M�B�h��Kn_��M�}2�3y�����> $ʕ�K��t���w9��j  ���D���AS�Z9ʇ�
3S�pG˯'갊"�EK<���[��D���т���N�I^�>7�=�|���:�����4�Q�&��N2U���ﺜ@�?p����R�h�J(T���|&O�_Ip�������H������U����:����v�����gW� �e)�=e�<��KC��v��9K��!�%�f�BRU���2g�2�_K��I\��tg�<�g3T���ӳqN@b1&S��F�q{�!O!�J��&�Q��`v�M�G��.�l%g�xfM��<�b�Οo2�Y%#��
�~�!�,���C�rO���+^;M���Г9F/ye�ML�xe%�9!���ڥr��vh�I�s:t��,n7������z��MhvG�	����)w��H�f����*�j; ��|,�=��g$�J#�EM�@eC��^��O�ږ�?`�O�C��刱����'�)���&4J�T Y�.b�n��Veb��������K���,Eց���SU�wp�$/H�2�V��el���)}��T���{o��\)�k�-(��<���+�����qE:
����$��hN �YI�,䆑B~s��*���?��OY5ͅb%XW��"H���}K�;r�#=9�vO�VP�p%UZ9o���N��� a��܃�*���u
����*5���6������`�⢯��ٙ�6�� �g]��&�N�t~D���4X��>L��=�/�6|��9��yɎ�����Ρз� �c�:��,0"����(�Q���^(������ϒ=-_Ғ3c�����Z��?j��~�ފ?W��������ͼU_������u���r�a�~8�$#�����|�Ta�!�Њĕ4�s��;~�s ���#�,{6v��q]@�� Chr0����t�Ϫ?������hF���ŵ��>V�C��_E�h^�H_�����j���%�;̏K���@�U!�ɔe� 4��өوu*��G���|��SHŎSݜToq�M���$�O`p�*ƥ��U�W���З�M����,�Z���`m�	5�;���rDCQq{
w�������j�2�z7�	� �O��Z�R����M��o�+���A��CN:�腺��@t��#Fn)%Z��YaT�[�>�؂��1�\�Y`���b��R}��L�g!�⊤�b�p:9a�^�fv���]Q���I��`��T�׆�`�y� �h�|8��P��@�ѻʭ9έ�Y�L��>!���\R7����������16�A�n���G��	��z����V?��`���0{e�b�<�i�¬����qD�~n��{D� ��ko�)��m�2���B�@�Bj����DY�+�׀9.�CYā�o�k�M�8 �� ��Z��Si��-i>V�J�wē�H�]��b�����)܈F�WI;g�Ay�贼�YpŴ�:�Y��cz��5�Cl-I{J�{m&���ö�;���bS�Ag�8�R|�I&�7��O�G��BdA���t��"WZ�0}��'W���S�lh6�)��+��!(
Q%:V�K�gJ�xp�������XF@r�j�n����c1�p�ƞ�?�9w�F�[c��+��H�@�b���2�O
��UqFL��,�aIaYm������&	s��<��t3;pڀy�����D���1�
W�kUR+(��hHIӉyIh������F�;E�dx�Lpn�4�����|�0�@DS��@�ZwY?�t���vf0����'��$���gci_��~g��L�����1�{��N�R ��w�+��d���Ϸ͑.'"���5voU.�1
���]��Д(�<�$��y�*���>�D-�?�n�@�`��d||�%�x�ό�J�S�-ٝ|�A�]�?/��ejj*:����]��p��=��NH���3je��A#F�8n7����G��gI l|k� b�/��[&p��u���7�G��Z>�LsTSN�,��0�j�Wv���I��V�z�Qp)С�si���|{������e ܎�sG�/Qhssm�@��B"�Cri�>��G�>z��뗟e-Q��TYь��;�W�$�E�� �fX?]��uM�2���Daa�8�Q�p�8���0��!e�I��r٥.[(ּX4�r�(�DT�غ�6�uK�|孳U
��Y��VT�g��Z��`�󸳰��i�[�e�O����QV�ۧ#�ٺ(4do�V�ɼ���G��5���]��{��qs�7鍳���¸�m
+R��ҍ��D3|}�z���1E 
�؏��w����=����2hn�j�m��(�|f.�i�&����e��!�-@C�e�\�uE��[G�5�F�f)�Q���
V�-�t�/xѢ}�@�rY1���Xt*����}��m�d��~
̕L:�?��t2'E���]�K�E�,[@%Nc��q.8�$h�|sɸ��ћ��_��h�HL,9K*Ϭ@#T
;�D��8�������+�\��_@w�:�En.:x�,tw��L-�\&��<���
R�nsh: 2�X�_"Ѥ�u{B܋yQ��<4�d�ig F:��z��ء�p@�00?m���1A��i� 0�PXlxV64EB    35ee     8d0XE6�=t��);�`����+��bm��E� ~�b���u&�~M6�WӤ���m0� ���{�\�.4WH���S�:z���B�G
���K����G��ׁ��AH�^K�H%J��eȾt!6���FZ�`0or'<h�1S�45��,R��r�8���6��u�V�5HE�{hKK�#ӯ�)�(�����;�~s�T06n�b�%�Z^I��/�i�e��]���g������ӌ�Oݰ��v��S��3�����6P#����e+KvԦ�s���fИ&�~�h����Uv-��n����A?����%k�he�:ܨ��&��*Wc��Z��û�r�anke��p�9K5�V�$�*�Z�����"�c�XU)��u}5<�	����@�ڀ9U�n݅5<��´H�~i�����Ik; �<���G�\՗]Z�$��D�'��i����}z�)HУ/�S��ty�1���0����|�"b/�2_�RZ�{�|w`�,;�@ƕ*+0M��MG/�h�A`���$�nU�]GV�,�����P�©����O�A߂s�n����s*�,��h[I<�n:�F��M��ē͵oL��?�FA��=�3�ர���[����<�0�|]�	[�MY~b��u����w��:y���Қs����?�5�6���"`5�Op�:�(�m��"����SR4r�֗�'���nA	��R�NISx�͊B�ݘ��)�ؾ>�d�.h��k��(�����o�؃�ԟ���{��@�en�˗� ��͜N�	������"�?QiA�=:۱b�g�oyr`CH��Ȧ+9+36"�\�����y l�2FYE��,)�E5���*�A4P�� ��ô/�����	�뒰�hy ��[a���3�jl�!�/�)�,)O%J�2ŧv�e�M����'x'~��0d�A�=�T�H�}O+�C�(9����s�����q�_��'.�ٽ�лM�lR��!��񣶐��$��#��O�K��B��e��d�[G	�쪷�J�_ �둚e[��C.�#���Y�3~��~F=b��~�fϨ�A���h�fk�����m1�/!f���Y'Ub�<C�
�B������m����O����벱ޗ
D��
�'���1'��	�@���Y�sIc���×�M�F��R#	�L}����x�cn-��O(uձZ��JEɫK���kx�;6����2��b�ͱʟ��3R��zzZN&�J����o���� �*�Σ}���n�H
�/��R��2̆��X7�0DG�~!�l���|�?��)���R�%N�]�6k���������ijĀ��L~�)��!P^L��~A���KJ�Y��3�C����EB��"J�l����.�[l�?�A����H
I�X>Q��
<�
m^���/���y\�.^V��IA;%���ε���P�,TE�!8��ਛ�'�i�\���?�e�e��� �>-�!�<�����2 E�1���i��fs�Э/�O���S���XZ����~O�e����1=\)Z.�h����ahn��i0�|��vh	�=dDk��O���4X�:�q�$�b��N�C����'�:�p�!;|����RHJ��ō�ޑH��ٕuS��;���g�+8<hm�5nF��͡U6��?�&wQ-\���"�v|����h���S'�S �����|	'[4�iG:;����9���hu]Rt~�Y��Ko�.C�%�������`��t���?���΢�_�����3�	��� }��*a��_��'������\23�޼_��+�4T}����h��N;���Zl:�S���=E`�W���n5&s�c�q�һ��g�ȱ=FN����&V'V%�{��O���).�;�S\`��(K�?�U� ���p��Ȟ�1��qA�Ӫ	����ۮ��*5�W}�1�e���F��y7�a�(�����4Ɗ�K�묰u4Ā�,g�=)ʦve �@yUD�Uq��S�>�˩������QdM��A�"�v���=���,�izO��̪��W�J}|�% �7�4O�ְ'��D�O���*YX���q߁�(;���s�#���z~rNg���:"��VET�E%>����x�_�6��a����M=�M�y'@��+xDYlL-��*-�>����0̑�1�NG�5p�vmi3�����0c�~0+�Κr�