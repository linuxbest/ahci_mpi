XlxV64EB    fa00    2f80 #��\�l�:���4�a5��O�k^[c5x���:	F��j
7��h�nB��%_�tD6��갧��#~HۀK��P^-��w��jXJ��+�A�뼯���%�c{�˹=o�3^��)�!q!A�Y28S@Z����v���p�j��Pv��
{����Z��_��f�,9YZe��R�C�l��,�>X�N�yKj%k|��*\�Eg�y���A��A�q}���>I�ܔ]f�4%'(2�J�c,WpFiw	�_�V����M�>�F����/no�������[����ު8���+�~^���������{]��R=	7�^P{L�a��U�P�Bv��F	I�ޡ��=Ɍa�e�wy������iI�W�����6]��L���g �+��}��O�XR�D��ʷY���lb�o��u0�nf�����f����?�V�Γp�dƤ`�C����!�X�C>�/�8�}�ɽ������Zp�������A�RH^3������۞|��r�^%'|���su��k]��du�T�lH�k/^i�Ak��93���w"3��cT��rk����d���ҽ��������p�+�.gN
� �+�Y}�p��6��
���C����Mz?��m$m����Z;l_�-.�? �	 �Hx#�|�J�B'ҍ$E~��(�$��OM3����-à�#�\����v1�tg_�������S�s�tk8P3��s�J��uYq�x�]���h��+�A�IO�`.耋�;���0YZ��X S����-�J�~U�����1F��R��0��Rq�@lT�"\β|v����kN��F����k䥘�m)~@Dk�������g<�Y,�0d��DW������Wl0U�R�=��Q� �/L2^i��Wh�yS<}����0���W�1��\���FQ���{<]t�ǤGq=w2����Ҷ'�w���u���R��/C��!�Fb��Cr�_������{�lq��t��$R� Ֆ�+.�Tj��?��T!�ư����w5W̷���������_
/���/g�+�'��b��>4�:��,p{msw5����!R%���o�NbyѼ�d���U@6���S�c��i�p\9_C]�m��h=����P8~[ftO��1��B�*�G��*�?F\Cp���0qr�{��D 0�f�z"�\�}wЪ�����ͷ>��5�˓�+����� }�RM$@4�ߞ!Q,hΝ�w&9���Iá�6��n��y��q�xy��o��[7.2�m*E8���Ӂ�)��N9w�Nƞ��c\X�.LG�����T�>!�%�ۜ8 ��#}�N�O�g�/�3]@
M}��MV߇��`(ʯo1��ƣ'@��o4�^�.�t�+h��<�3����S3�dh��H��I�!~�RUu�[��bM�U�ۆ���U(M�|U�3Ui��@��A8�ޅ��5����9��@zMԂ�; ���;}�ţ2~���K�h�@�d�?�O�NL�0�0G"�6���s1���0q�ǎp�&��\D'%���ޠ�.N|`����զ�L�[r� ޯ�6��2W��."#�@���LDk�E�F���f��ָ��b��9E�Ìh��sAZn�6��m�`�c����>�g��	6�I�̌ۅ�\ f����U�dђ��}(�݌h�J�  �$ѯ�+��#~�:�|C'�c��Iw�M��	<y��R�%��PMG��\+9K�5�T&N!��;����N�d�Ÿ���ҭ��$�?�}�{��>{u<Q�9�C�s(�@��j&ܳ͠u�1n�7�q_[rw#=�=��,�.�����1;��?Bw杺BX��frQ0�o�/p�7&�4�c�R��-*R8�f���A��acH���
�a0NG]p���m��	��휞ˌ�S_�aMj�:A���(Ɨ-��Ϥv�k-27���e���&�{!^�b�䙵�Hv�
(^��@���ҍක�d	��X���tZ���X��H7+�g�nxn4g��ɉ#��Gr<�CG��%5���H�J���R��X���V��x/�ɧ�Sl4.B��{��
�ֆ�y�q6h��~���uk�"���۾�N�^)��vO����a�bC�R���ϸ���Wi�|<_Q��.�712�rخH��^�j���

�Lq��h9���wLS"sX��?�̂��\�B\�[�ա���d�����q��єX���δ[�-
V��w�y�Q/*�mRb}|��$#�F&�G�f2����h��̃�=�F�NM��j��V/U���ۻ&�;yb���50��BJ"r��1������a�%AҶ�`]z�т�	@������F����{/���#u�jI�=>5�^7��ʊ8|gw�%�~�f*̿�6�`���J�3��4eIv����m�O���S��.�aђN����S�R��MN�g�6�A��F#l�Ǳ��[;a��wދ�J���u�>�@T�J�$����QR���I7�|׍vA8�B���Fr2Ђ����MQܯ2w�bt�0��rEEK�o9����b��Z�`<��Xho+ےU��Ǖ%�5~�~+(�p���G�#|�4(/iiG�n8A�r���2�f�4eR�)���f)��[^-T`�����`~Z��<�@#>�7!8Ԡ��ϲ?�)��~X��dI�Yr�ƲĦV@`�{*��9�ۤ��h�ʏsdT3�u����B�� S��&���M�Z�%����^��\�fU�:�ճ�K��:�"m�q�Fq$%X�4b�^k�;�D��;5�j�8�,v�?U&��XC�a�o>��'�Z�C?V������&��j�����ٙ>ߒfA�'7[_m�o��'A���O�����;*���\�3je(ȷ��yFE���/?D���b,��g8ہOt{i�#={q�¸�_@�8!�rN�}	>5�\x�	l.ƀ�#J����j�}�0W���YW�KN��g�Z:BC=L�ߨ 8}Hۀ��I���z#|��K�1%����rP���	�ܭ����3��<@t�m�L�kMx\�gr���P���P]�=�����eae�x��Eв�!{��[�rӼ�$�N޼�/bm��E����6w�b`���/��2�j�U̕�vι;�ѳȋd�CKQ���!8��N���v#Mi���^�;��{9/%�)>�sC���Y:����*Y܈F~��x1͏�AX*�V�K�d ,)�rl�m�{�ݯ�����d���70a+��1�y��ߨ:��S#�Uų�*��	U!Ԫ���֥����s��i���qv�YƐ��%k�0�\;�G#n��Ke����?zmZ'pe7zܞ��%u�n<"j}�2�YU��~�){!����Π�掋�c¥�k���eֱ�8�d�ܼLO��͓�U�~"�a�_NR�Dq
.�U;��[�C��j�3��43���&�P�֧n���&V�6�Z}�HE=�9g���B��ێ@����~?.�1��Z�o04�2��$Ĉ�JA��~�o�p�)�0����%:���sN��l���<���#YhB��Eq���EI�qH`S�;\.�Nw!�w�c��1�(���B�E_�PnH����1Z���O��X�A��ׇ��[�ܾ+tڴ���Ӓ]�C�y�(>��mc-����r��W,߮(v�
=S*�,��yl[�"I>�ϝ��A!,��x�M�.4|�͉�8-�t�� /�0�����߻X��n�� ^(o9��bJD,�`�y���p���@w^޺��p�]<�GYP��G��u���ψ��X���,ϕ�5����[��2M�eG�W��8��?�T
��3ZKX�~�	J(��;%njK�e�׈�G��g�z��'��ےJSmP�֜X��K0���ಈ���^����A�.%V�Ş}V�4k����u��9 ������E�+W�=)_E�g<�w�G�g�k�W3/Q�b?��h0�nD�>����L�E*�Y�.�nN��y��D���e�����,�W�9`��Q�n�Y��a���@)��?y��(��Sխ�^���f_��;r���(��v��/�F�E���� �b�Q���
��W�J*�y2���y��\쳏C��m�U�l.�i" ����䱋+�9�gFy7��3p�/�������`";��v�Ֆi1dq��8R>C��+=@#�Q��Ys*�Y���o�Bt�ݴ���kLfj�aX�Q�L��'��$���6=��o�'S'�Y"7w���L?�oEgY8�(f+��]#���o�s<Hћ J5����d�/Y* ?Ѕ�h×�Pߒ����Df]��P��-�?&�'��f��<���W�LT�Y�7hO�"��|DH
��ꊌ�G�D�?�G��
M܆����*QN��R�6A��e[hW{nv^wP�	b�w���P�(���Q�K;��c؃�򷯅��6�����q�J���N��W�Æ���	U�!|�H�^��,�(.�J�� � E���?��f=�R�]��A������~,��qe���U|h�U����j�ƍ� ���.Oc(�#Qdל#7#��@�����E;��"	�[�Θ5P�n|��7(�X�{��Ձ����!j�JQrP`|M�+K�a���橈X�T4D/�8�^����J�(4\>h�֚8�	�@҂;u�`���֪$�.G4�Mou�	!whM��jY�>{��;��ǚO_��A�U	C��9���}�鈚����2�9�㤴c����SĎ�x�c��sIZ���o��}`�������:��;��Y+�R���3H���氟�$��͖Cn�P���$�n�`KtFp�!���/�O�dkt�8K�JM�-�[��O~����o��pu�����6"*�3
7RT'�X��b�Q7N-�ĈY�VFJ�����������~f���ߣ�����,U�a��i`-�6Hu
ȵK���g���N��L��4�HUE/`S>��N�)I�m9��ќ��ɂ_i;�MÍ?�L�2�6ϋ5vS��!Ǥ#uN2��	����l�f�5G�<��*bc�`��l��pL��Sٖނ����~�_�K�� �N"眹�7K:�͸0ix�<v���������n�/��5M|I&WUk����uKƮ�j���)����?1��c���/fѠ*U|pƜj�\d����ug^���R>��2�/�����E]�����Fr�ܭ>k��K&ϊ�	p�h�����-�p�d=�0Iu�ġ�T�Y�݅�h�sҙ3�k��KYM�����3ث��A$5ۯ_�-����f�D��H�7�1j2yeU���|?v�]��7�Dj��d��Nz�N�~}�R,ĄR6Z�m�1�K���n�����-��:�)����=rls��������c6N��4Ғ-m>_홚�k��u!�����"+�f�w�i.˜��qE �zp@���H�����;�/0��=Ad�΄?�̅��; � �8Rdp�UlZ����~Wva���M0�-����f����y�G�*�'X�������F���-ۮ���ٽE
���L�t�]0o 9n�C��c��~sj��/�BA��ح�ǟu�J)R�TG`n!�89w�6�h���r�s�7Jk��@��\���XfmiX��͂T{������v*�<[�
�5�Xg��3OjԲUl�ZB��Dzy���<&���y��f�0źa(Y�G�j}{5�ϲ'�]x|�3��/��A���V��1մ:�+1��"�x��sH6�����:#�GX~Y��n�D�u� G�2Ĳm�ء�e#~e4��a��4��<a[�'�ۑ�4&`x���W��ꐢ��l�ZI�A�]@o��FZ�!ko�w(@�Eag���ƀ۝�U��*��Ud��|���2�~=�z��Cl441�|���bn�c�[X��������^R�H�Pa��I'�R���ooo�� �n	����^`�]�W��������l��*a'�봔4S��P�"��y�\��?q�y�#��	�\�W�f��&|Lx��L��>D<A�t2%��|�K��?�rO���Z}G�4����j0�c����#����k�)���Gv
�7�����A�\6�̛z
�X�K�UC�#ĲE�z��~�A*B���׃	/�+=Q����}�j<R�O./>� T�Wfevd��|��k��H�z��J00���(x�X�]941��yq�I]����\�oB�#]7�=$��g4��dd�Mx2�1�gw.��v}��P[�S�n��%��A�d�"#��o|*R+.'�ϫ�ޓ_����J_0��x�� 2��wM�h�U;h4���t.ҧ�;��@P�o����䀔4��~�X�\�����p����S'�r���9��Dw�� ��8=�Bz�� � 	y�&CXq�

���qM��-1C��z�J��}�,��?�u�%n���b�U���*�nHWf��4]:8$vƱNT��6v0ok5�;J?��OO�M��׽˃�g
I� ����M�P�%��`�T��wX�F^i���E��R�WS��ɳ��ӎ��"�I�&(�,ީ�?���u�M[�Kկ0��:r��Q�cY�[W�7�o�D��4ֺNI[�cs�7��;&|-n�˕�~���	�2�?}F�፹S�D��i��#|	 �[���	,��zHX�������,�����(i��!�E����#�tԋ�{�Ʉ8�'���&4*ѻ�)ӿ�9l©_Y"����q��I���w������twN��g���z��0�Orf~�Q��3Xg�Do��޲@��/o�; 5+���Mp�s�Q8�1Z|+.�{���1�6)p=L� ������e S�����������b�����!{�Y��7FTt�Iz�!��d+)%��=IH8 ���b_L^8x��(��S �v˶ts����[�[$����5I�`���g��rc����j�pj�G�SL"��N�}�`U�����K�mV��M�V8�J������>�*^�;$3��U�A [W��|3�x�_'K )��sǵ�(ѿ=�aS�Yp��9r�(u�F�S��D�>櫱��ʅ�l#�}K��C�&�]�z���{䓋�Zcj{��4k��9�Q���U�
�Vad�HU�Ş�ȃ���Nծ kbuZ~Yv��WHH��y�¹�3�~ =��4��� w̋x�S����/4��W�c�Q"]���-M,��j�VI�Rm�=eG$c��U0o-C˗(�D�X��_g޼&D�K#�	�=C���b������b�T3n�{�sPH��;�42��QϏ�ح�naӌդ]�� ���Z)�ȀYS]b]b�n�4�����3bfwef6�˨��J��gM�-RQ�v�e�\\�(�Y�)�hm�6�DP���S��}[Gh7�SZ��Zs-^��	��i�v�6�����-5���&��L�1.�������N���{첥b���T������Bv_D���0~R����Yg���g��o�-n���J�s;j^ v?���8���=�	�Q��W*��C�Q]I�rI�YA d&�����E
��s����%�M@�;m��;k�4?�VM����%�R��C!Օ"2�ǚ��39�~kx��a�oB�(*x�)p��ȯv��G?��ITϾ���A�U\�3�� ��Na<�H�KT�g5����t?�t��y!��N(8	?�i��@�2�ٕi�t�(�Ӭf���>{cƈb��L�YY��C�sfO�HKV����7L'b'H��M,�5D�'��Q�N)�~ᗈ�b}�fH�����z,�C-\-�VR�#F�[kD�S���Gn$�.�.݂�4�^�ۆ�<G�Nt��d�Bp"d��ba������H�h����r�v3s�֙�NR�{L�";����{Z�o4��]FϷ,���������8�llt�)��?�,\����Y'�eyE�	�Z`Ci���tO
4#qx��w6N�pH�H`bzC��,����O6q���(ݏ+�饔b_�����dJ�~����c�>�5�L�r�@Ջt1$Zd	y��<�1�0RQ'*�0�q/��+C�}����VN����%>1[��
<�X?���}�0f�@�Q�`�����LD���J�+%���p4�f��Z���i���1b��V~~9g���#��]�#:[h���v�p���{'�P�χ�B�/\xP��Z_\����;��N���Z�g��C�����7OR?�f�NuZc鬼^�F�Z�'�h��oE��a9�Ѡ:�5[�ٷp�.JU'�nn�7��d>�	P�ñ٥E� �@�=;f~�&ImD�j��.��*� ���!
��'�U�E���Oq���ŋ=ˀ<�`��&h���z��|5�qZ��-��d�����<����[����
�Z��i�八���|���_�������0���o�be�}�^M����'�5��v�MF0��<������G�ؖvI�GJ�x�~ft�"f�w��@�`�'KV���\U��s3ײ�-O�O�t�9��cq�C-V�k�_#���uB-Y�Z:>��>� �p�K��.�J}�@�S����H��pP:b�Q��9�����'U�0��_����9]��
�O^q����[�o�1�Ѥf`H�Q<| ��[�U�j���c�9�H͎O,Ea�����E�`���O�=�9/3�Ve?ݙ�Ɯ�\FEe���Gsq�bHe!�
y�ϰ>�*�'�՚@5ۙJSl��lH''p����޲|�2
�"P&Қ�����c��ҩT{e(y���;@άl���l�'�#(��W��ګ�1I���N�yR�R�I]5�F�����E��.�X1�Ll�N��H�2ͳ���b�{7���7C�r$ Q���]����ߑ���,�rQw���6\X[��}��:�-�;���!��*iL��13���5T9�|X(F��<�Y�EE�ׂX<6c-X����Ϸ����P�>>Z��<G��Q�ι�d�SZ�-?`�̜��5�c�i�y������[��������������_o)A�jvq� {P�<Ԑ�i�N��9�X��/2+���O)���K��Ot�]��ר��UNb?F�#m��Q�4�~�^}���m����A3u=��N�x�ϝ���k�"�o�����n��\{��:CK�w���vڊ��}�N�]D5<{���=���OS
��Ћ׿m�V��5�k�H���^R���O��R�O���&O���}�E����A�]�W�a4�-�V�DL"�	��<�Ttƿp&6�T;��8�c'�mub�*9�NT����@�8�߿Sd��N��OHR��5��Q�{8�	0�>��ǜ��7�g5����t��b���!��z��h.?J)\m�i�s��-I���Wa
0�.��Y5{ �9�#���50u�Nj����g�4���¼ ���ҫ�	ʫ�38>�XY�	�͝�k-P wA���8�C�t�G%
2�9�s��`���<�g�}�y�OJ�ݢc��:�Pa��+@��$�s�7q�g���½5Uq��x:����06bh��������^Ӂ���ޮ֠:y*�^��)��FS��*�@�����
����傼ٖ�ti�?�[	���x��U�?���,�(���l�>����׼N�]_�f�1�j����[�?��Xg6R6?Ld��TV鯼��~� ��"�PF��Ni����I��(��\pUa�P�����
��dXp���\���i���`�+�:�}���h�.�dSRDm?�iH�t�ѽ1�;J���yA/
�Ӽ���SK�=��f���ttͧ?_�������W�.��F�KiY/1���+��}�;���b$��}� �2��onj���}zX��A2��E�=�-_6��E�Y�pY�c���>c����pZ,�R�1;b$6��0��sV}��n>��H��vT�@�Db�1��1��8�Kզ0dJ���( UC�T�{��x��	v$�wd���C���?7�aż��Yh��e�o����O�s��������g��&=b����2O�_ו�ބMp+с��7��J--J�21*�B�d�v�{͑�j�14��*��|�7-��W�i�Vu�p�tf=O/r��E#���N8R|��6nr���ti�g_�ʘ��TqO�S9к���~B��cnn!��a�5͞d-ѽ��E�U_ذ?
�\��Je~�0͠�UJTċ�g�%���,��"�!;��Bm�
�z��N�B:k���CS�ͺY��x�d���Ayr+x%F2�MFQ���c$������0�G�:�|R�������SC�����e,9qˢ߇NT�Ǫ?��ă�L��,���_p��D�>�sJ��)<+~�B��:�0�8=60:w>��^��voLbR�?�
G1�"�[��"|�6�9��(��I=��aT'��:�έ>�A���w����8y��ԙXR���&���?G���g�zg�[��\y��h����Lo�I烥�Ζt���7Z�"���uQ���f����(�����7gU{�/:�F?�?��G��ޮ���i�pp��W�Cxg�>j��|͞�ܑn�H�͖4uw���ʪ2��+tt���t.�(�7gnp����$,�yaD��iW�#��+���ͭK�;��W�W��i��~侒�����/:��j�m��
S$���P[Xǫ	���ۗV���F`CuA�rI�3J2G[��._�7�-�Q�]�<�aP��d��F�y�IQ�+�cw��D=z��?]u��5dě ����M��n�0�T&�(&_|�3ޟu&S��\� Mp��奁�\ը���S����߭jY�*$���J�?o
������@�[��kKn��� 馶S	õ'����D���5/��[=Z�@�Ɓ+P{��m���	�AvPt���1�̨.�-פ����C��]�^yѽؙ)��5� �2��VGo_���[g�0�A���ꢘc=eHȠu_u�\_SVR�eR�
�b�}	Ŝ�A)'���8��b"7����Gh}�sUV5�Z�>����r���U�1��_euk���g��?�2,2h"�sV���I��n1�����9�^�{3Jv�<��*X<�F�]. 9a��7c�j�d�R�C��a��y�+�H�ɋ�d�B(G^>����e���Q^�KL����ВL��E�B��)��>z��S!5�(^l͙-W�5	X��@�LA;�I!۽uěcd�� R�]g%�#w��^5o��t���a)���׹d%�ü4��+���fx�}1'�uv�*gP�����R�]�SQ�fMx<R	0<���-?���O�X�ޱ�}���*�U9����5��ꥨ�[�c�%u���A�?�"E`�akH����K�mms�l즳�vD\������z�
w$�'j���f���_��R��&c2�C^�s��%�Z����d�*��A�\A�g9Ky�6�"q��>��w2� ]J�E	�I�	��M�!�tbߐ?GE;*A+��䢖^��g��p�q;�˾a�[�/:������W� �"�N�q"[%��g�	�g�n���o`/�v��zc(w%Ä|����g+���(4�G��d��L��7N�~'��H�~�1Y��A�I-�[,�^�����̀���ro�2�swP��V{�J�g�}U̮�s��,$
���J-9�b+��\}�[J�A����\`�Q���#��ޕu8�O;?
WY`�rL�Z1�4�V��k)�uEHGJ�����*\U�zaY&�ᮃ��ԅ����dm���K(��En���+W+v �� ������T%���'ZO{ѡ��Ve@2Ł����?'��0��4	EWM&�F��;	�=�ܲ{��k�����/{�#�8�� -m΅����8��T\(uv�z�pf ؖJ/e�,i��s7�ú��,�����;
��7��2�XlxV64EB    fa00    2a80,Z�begPhv�I`n��$B|��γ����;�u���=��,4��"��J��C����	�k8%��X�|�Ԋ�i�M��4��<!z��@�����H>�<�(�;M���4#v��3q;ۻTXn�#�s�,`�b���,<'�nN	8Z�����W{�ұ���z��z}+l����nCQ����@ ��ѣ��Rf��!*���e��Dfz竼�k���@98�"[���i���zE�rndFz���_�C��lH�J�V:�D|m�v:߯-����M)���8�(�cx�)֚�7���7�g8�F�I�^憜��n5⺿d�xT�
�9�O@�׹�~����XP<�'+�֠T��ǋ�����&�r6q:�sw���!@K�e����(�����vH���HQ˾>�p�_�:��T݌��Δ�E�܃��?��W�ST�[�=��ggE'�r*�0��VvIČ8�L��w&I�x��R� 
��R�@��[�%c}��N�j��3����B�{'El� �W.��CX��l��u\a4B�;�r�z�"�fBi���91�b5�O�1ū5�y4��;ƭ�L�0��{7����D����;��3��Mf!���.�6Hڿ�}(����<!�N�СC�n`�C}�fa�{f���"y.��?���������M@�l��	a�`��㍠���K�+@�Y�`˘(C�x��(�݇e�l�����}��@�;�p�^��U�4\R`�C���"b���$D'�\��B�:Ca��d�B��i?,�J�}��L������ϫ�6���CX�����jS 볥�<1��Zh���U�+~g����A(���*��ְ�Iѹ�3��5)]Ԓy�س$���kd�24Q�G>-��V�
)t=>���&Z����/�`1�Q��P��Ŀ����� ��01Zshn/OzD*�X�5Q��$@N����ldQ(�B��b�=~�Υ��8�n�h�L����<�%�·�g����3��	�<�l!��8*U��t�m�W�i�<�+���䤀�%�$�\((�0
K�Xޯ��!/�C�n��-U)eR�,e��j��F�.�I>'�]A��W��n�����p�b��2E����u`:���7�+��i�(E��	�/�sN��v��a��j�r:��W!�zK ��F�8f��+�ΛL���6=U��_`�����rj�[yC��Q�̾��{R��WMvd`�KeD�mZ�v��D�i����q!� ��2�k��	|��K�����Nr�l�]������i�j��*/��:Vp,S׈��I~����V�I���U��%�?6��'o�{*UC<١r'.�9��m)�6�|����9�XqkE����(X�����~�7s�f���&���*$�!z��t0+����hx�ڍ/gl��0�%Zv(�.JG�gv���4A������������د�.C2��[?������(��ސ�,2��H�1�c�9kY B��<Q�����J�ғ�^��m=G����a����t�F7s��`�F�W�}���j��ubj�+0Uy��Jh���p�+Q�~IP��2U�I���$(�η��;
�p�8׊�9��S�4�} f�P5Ξ�*���r9l��^4n��Lʽ�u0��5�������G���YE
b�d2�Q:���ě�k�%���ō��7��>F�T����v���#��2,���K����T�w���1�@����K�H�T%��$m�=4p�o�<�*�r�ܽM��Ѵ.ﳖ	�~��h��u��X�_KT�����	18���c�
�m���u����A���l�O;2{XJ�X�^�?���d�EH�N!�׭��	���=��Px�-A��z%�1��J	#�
�&*.�-���N�I�$��"r~J��!�ms�v\��'6�a�����j�>)����8�F"R��$%�p����c@�y��M
���P" ������?�PX��]孳�E��9'd��\����8��R�v\DJ�D+B��
0��d���Һ?ZJ7����^�'�#�7,w��5��[>��R���`���`��w�gD�텸<��T�/!���x���ܕ p8�f�6������
Y'�8�_�!̙���u�f ) �S��*#go28H152W�_EߋϧE6-ç��?����t��3v�$�`�����fN���P7ڢ5F��禹/4 ���߿�Sa�[�����5�.-�C����n0�	>���ֱ�a�,���($�9���&�u����(S�	�����Y�U?�"��ҩy���n�!��Y�<���&DW�2U��8��o�ӥ�*�e?��-���&~[9 Mȉ��C��@�8�O2�0ޕ5O��a^;���|�B�k���-��\O,���ʎ��wء������)��%ϯ���SU�����x{%�i״��"�b��䋌!�/�)`[[#�c(˶�10�b�<B��[��o���M���C*>����^���)�빶*����>�6�,+߾�R�Q=� ��;ۯ���z��gr�;H�����qa<�We��k�S�����36���oFMJj=-jl�����PoG�v��&)�h6�W�V,
{`��\Aȿ���ڋ�������Y��qH���-�\'���Q'8�`�G�S�f��(F~6_�:r5�Z!��۫�k�u��x�ē'w�9,�Exť�`��nd�O��'���
�+֨�R�%�5Ad���{T.-�RJ�T�������%�L=�(�p�Z���ۿ�<��e&h���U��%,��6���Vd��y����*� pҚybn�܇^��VQr@X���>֢1��5J���*�:;�?�T��h�jU]P��=�d2A�`�{v�*�\Y�*
F�;�tHh`���>j��&����8��)89فt��x�<zV�s�j*��o�ǐ�Q>o��B���S�6�rev��Г�}%T}}���7 �:m�)���Uc����mŭ���E��9>;Y'j�~v�k_PР��X�c	C^�1�6{�"�Ǥ�[�҇��D/����#LfŶ�*�C�-9霤-�<�Ӌ�cw��+g�_�'�d�I�>wk�$	�L)g-}����}5h�d��"Y�&��1݄��y�*�aY�WB��	�ߝ���1����1wXV��r�p��S W�#M(���0]Y�.\��Ŭ��/�����}��.�� �U2G ��%ﲸU�l��k /��!Y\���u�@U�$�^'�J{�ݔXA�8p�6T��'m��q沐�u������QzM�6Z �-��* ���٧�>��z�����ti΃D���G&�S�x�Z5�V�$%yG:s[��ZY�¯^k��U	�L�8>�.�ᙻǴ�&X��|pJ,��]Ŝ��#~!N�C����Rz�S�-��@i�����5�J�*�W��x��󛹜X��#���,?Y�b$���O홛|�����~�����n�����_ģ�K#�"%#�z�Q㥶Dr\U�Rb̑O��`76����Ⱦ_;w�~E�b�A��Yvhd��/��þ������؊!�vT�gk�(��s�D��uΊ�>��VMa=A'�$�~s{���������x`����.U������#��4w�k�t���?p9��e���+���c&��=	>��!�똢���	p:����l�,��F(sW�r���s���S��%�g+~kyX��T���ˣ�⫓2�ǳ�a3�޴V�����RY���W����#F8*����X��r�>�6�I*�bo�6���͚�� م�Ϻ�����j�~���gsNȠ�w{>�5#���ǥ�&n~PI��4���n�Czʎ�o������Ʃ�A�F���	�2!���oF���0�PK�k�Xwē�&������	s}T�T��!��|o9|9l����47\G����" ������g2���>�{��ˤ�{l�K"��s���Pm�u���������l+�s,�{��ss�㙓{��+[�O[;p9ɺ��&�O�e?�',�c��zu�#f �1�ԃ8���_2BD�ܫ�i�Ӄ�S6�8��Z��
a{���$�� �"IP���\F�zW�6�ֆv1P��{��5bʃ��-�|[=��bx��}+%z+�"�2u_`��s�U౱Lz�2��U��F����yK�9xH^�_|�ɍo���'�����g�V�>na	aאĺ���������-W��ĳ��&�^���%s�7�"r!��?�^��Նz��+ڵHp�Z�9���LE��ݟn�����d˘�6��c�ߨ�u�ġE�96,�9v�dl:p��*E4!O>[Nt�b��s�.I��"�����]M�cY�޳x/_g\ƺ�)�X!��f���^�0��Ih���l���O��l�#�w�d_1��O!���TI!ӋL�i�h���� �c ���q�(��,c�0G`�����ox�[B��ɀ��n���f�����]��Z�I��|����$6��I��V���&�y'5�H��������,(�s�	�$B|B�ՅT�{ A�(��mѺYE�q�ή�3�Q��З�����2ZÐ�/u/w�b��ܔs�CS�g�X��C�9��z�j�\�:蹇�l�Y�#�!�����/�YƠ�~�VHZ�&R�K�>7��h&�{w@Id8偲���k�zu����ÄntC�HG���ś���4�3ք�ehؙ������ޔ�k.�;��W(�K ������A�##�#U��:��Ů���BB���&������Lw�b�r�MHT��}�A`�/�p�zr�r����u��3&��s��́O� ��T�;��ga�`�}t��M��6	i��3��"�I���Ď��,+n~�u=g'�ѱ�HR��{n3?ca����՝��8hd[M�𗻆H��~���7
��U("�̴�a	M��t�0������_�s3�&���F��=؇|�ׄg��h�/�\�R3W'=֩�䝒n��86�"����ʚ����jO_�y.鍢���m�$`�)��6��m�4d��!=�8��+sx|"��~e�HC�#�,>2�;��a�K[�%�����ދl�s���):lE�8���(Iӱߔ*Bh���kb����.����4��J�w��}(3�u4�@��P0�ڛ���\vٹ�^�A[���]I{���_$��rA�a���w�&H�G�y�|���y#M�-�q@h� ��Я}�������=.8�_Ϸr�~��f��⟩�s�d���Q�V>���X��ЕdA�U��c���+�A�������eq�=�.4�PuD~}e�;J�ַ�K�$Vl���!y���9|��gG��W��w+�n�ۨ�j1�B>p�~_4oGʫv��ֶ��r���u�~��R&�|YLU�q�C��F@c��|���!�CTi;X&L��4��t�#W�ϋ9�Ib�j����]c>+��*?�ʴ�y�ًm����c
g �A�	�1`Z�:�4zc2yU?�v��6O�C����l��u4���AAm���S�q� �W�~jv�N:�´��f4
�)5��[q���6���k>�]YXw��(F�S�����T��K�{t�8�o��~���l��~����6o?��>��A�ZQ�ˮ����|q���ɓ�8'�:=>}iE*�� �M'��Iw:��y���+5�����/wҨܮw��)(�R�t)S�c;"�>��+bs	<|��?���l���������G�^nf![�����m�
��>O6W�{F�u�/!������Q4��焉�C�� ȤM��ЃC]'�eӭr�M ��:��9�����H���fs������:�jxf�8mx��؃5#���T���4e���c��q\�\�Wc�B.�)7e�$ԋ��Bl�Ċ�E�l-D����:���`2#�Z��d�9:�S+C��« X��70<8𖳛
~urC>o�rv��'FD��w�B��n����+>��_���2M:s��ˬ���
̆tp�%˚\{��fM�Eݰ@����: R�4�̌t�py��pQ���_D�f{#�~v]r��n �=�oF?���W/1	��;�~����ӌ^��(�:����aJ�e�?�2u��H���1��Y,���?�p�!�����Ab�WM	�;��X	�w��p����.�.,~Va�_l�]�+��(>�&�����'�D��T!���2�ܛ������/T3��ˎ�	��] E�ŷ�@z[���P�2��T"�R��x���=~޵=fq��n�)~8�nN'�Xji�7��Wpu��;5�� �+1 l�6���!�T�O/F�A��o�y�>���jD4n�K/�����P��1� ��4>��)@�v9;�gM��y��w��Ҝ��׀Ż��Kzݵ��b��C��H�������*jR%l�������jP
�Fh�ŷSJ �[����������Id�Tjt����:ʽߩ{&/�"=��'ݖ�j ٛἇLg����^�t���{�L��ӑ�=��>�7s�E]�6�]�{����]KՆ�Sgn{^F��hkU��P�`,��OЙZ�f��$G� Enާ��˯���̑�g	#�U��	��T
9yv��ǈ�/���aJ7A���g@��}� ���KK��-�{攓^f�^��k��-�����v�2'����ӜYY|����\�.���삮tu�(u!ᵷ>[������U��+��/��'[�5��&U°e���6ѭ'��3;6��v�!..�������gZ�؜kQ��j�%kDCp��sڌ����el���Cu
sW��1b�4|�N&a|j�2�|���)%:��J�evK�tm�,��B������V����0�ɿ���?+A�@|Y,.g��d�yȇ��w�x�e�	!��ζF��h<�y�šF�U�9O��|��_A�^��7�q�X���>�w�ډ[�����y9Wy�|��=\���UE�T��KgH�ߚ��瀋���ޏj�n��12K�򫚏�t����l�%��P�J8�ʌ�����X�k�g��g����U�X���A>��N��r~�;��f�#��%���S�����*��m-�N��V��}b�L� 5
0�B����Ѧ%�/���U���� -��+P;Y'B��a~^�0�F8�iV?HһT_`V����J�\�'��T��;���/���9�}L���M���E��-"��d�1ᓌ��S�(�Z��@�@;��߼�#�0��XYhp���Z�� �(?�Y+�����
�>)r�R^H�/\��^d���=7S�I+���qⳖ��#�_��rz��0�0�X��}WϾ
c��AT�bzP�?�2�!�����=�l�T�JO�	��L�;�2��9+5H�<�:0G6�x�Wx�mc)�V���W��ꔡ�zE�3&�MM�h1�8�B+�!.�8�[A�7[h�4v��ng#�D�2	��2�P�����'��]N�ˋ��ټ���Uk�A/tx|�S߭�|�V�x�I�)�_��DOS[#��#���7�"�-8�V?	��n�-�8�o�A9���߱�>�K-fs��O��� �O��mE��b�ɦ�q�]?
�?6�G�`k���o��"ҕ��IlM��� PӨ٠�_�AE ����W�ؠ�pK�62��L[�$��۫֠�݅��">w���
X��f�N�Qc��H��=�W��A�Op)�W��3kq��g�6���OL��>���d$���)X<U��he��t2~�g]��o���~;ˈ�y������3a��+�t���M�$o�OK�>�Ԟok��*������B��#�^��>D?�A��@V������	E�?8n��-f�[a���2�:C�8/9I�??411�G�Dly��"�4�[�:��1��z�=]gŹuFI~BәA程�l��P��{��Q��w�oקs,`QܕP��3��	ͅrY
6� �Lķ�2a�91��U�w��KoQg��;�EC�B��ۿ��\��#nG��{L�H.�P����qu�2�uiB�a��ٔ��ڢuk�K�~����{)�����"�(�1�R�{�B��]D�$�<ᣛ�aG�q�����S�}�0u' �Mq��J2���s����] �)��n�_��;�)��N�".�[������߮P.y�	.�_�D�ݸ��<l�"���%���g�rŲ��s�;,�st�f�|"�y*Mk�;A��,t1�����^m�dkQm� �u�T��tj��8Z�_�8�e$�KS H盔+�����މكqy��a�_��A%Y�c�]fj�฾xx>���f�f]EjM�c�B�  ��DK�VҤ�,�z��JM�R̢�Z1*�cfie��b1C@3����l�{[�U�3�k	��,��Pd��wvJB�w�Q�yu�9��9��#8�j_�7z��3���zOM%��n����I4��An���Z\�%v�E��\<��Y>�/
̤��D�h�vP;n��ky�8����
f�OyW��
��H�J��줪�X&	�	�Jo��ڃĈjq�Y��W�ec5��ƌ���n�S;f�K�@W��8�L��V������QO�H�O���hh�X<hw�|Wà���7a�U]G 쐀_��Z����]%�@z�GF�rO0D�W�Bk���x�<߹����vԡ��-���r��e$�웷�S�v��{$�ɢQ��}�\�r͂�'���zX��뇟����M�ش��WUE�U��@�����P�{npi�(�}�Ұ���xjm�	��w�Nဃ���&'��,�J����(ϟC���yQ�5B�]��VH���O�й�g�'~q�*N�T����O���^��� Z&4Κ!��b���B��x��Ń9�qS<��iB�Y�
��mh�\�.�8�ͥB�8�.��Էu~��־z����ý��HP�X��$�@��Nhj/=���x��BGk��C��X��O���:E�^�We��a��v��.X�/U�n��?ـ�%m������)Pk�G�{?��kQ�#s#��X��%���@�EY��ۥ/+��6+�HI��s����z���l0�E���o~b����))w^h�o'��D�P$D��P�����%β�/o�,���L�x�b~�Ց�ϼXK[f���Q��+HQ9�݉�|�������e��8�.�}���tB�B���T�Щ-6�di��]�F#L�0ͤ�n�i�V߃��4,c�ݯ�9/�v5da�*b��CʍSXȽ�L�;��Z�)Ͱ�@7	�~��1����E�hL�^�^��p�~b�b͟�ҵ�Hɴ�-�W���¼ 	P�Ў�k�4f�� K��f�����$���Btb>��U���O�FS@U���z�|�=kL��H�G�$����i$we�[.:���@��3T�A�z�����%�m�����f��o�KM1Vc/�@�ރ��N�� ~�3u$�Bc��/G@	k9_xtޗ�q��1��博܄�b�Աu*�Mu��+�A!`g�?8���_�D���l��]����.��җ��1�&uͫz	�nݖ໻�r�>�?����T�h�1����S�Ex�acoL�c	m�u��mE��S�v���ݩd�U{ɶt?+ ��=���TFIny�md���+�7�>�"��Mt�L�>[6�4�,�3�7��D@��8j����0ǘB������6'�fE���@��0c=������@T�&���E-3񚰵���;������Ӎr�'�s�}$o[�1��qd��z �}u�G��3���(-k�Q�"DMjK�@��L}�`�!@�?���=��P��Sň�J��}�f��{N��$�(N;��BPQ�Si+|4�,
���
E.�G���Ӗ�o���(<6�v4}Q���������l�n,�4Hb�5Q��N�w��@�Y��Oə�+kJ��1�> �i�n�o�T�B��
�d��/s^X��,���1j��cA�=v ݿ�8�&80CS�{g�@:ԑe�5�ĸO�(_�8�X�=0m�o�i%�Ft���D�5$`�R��KTK׬+Z�Z 鉗:H|�L0Ŗj��>���H����Mp��Ǎ{���f����xud�֢j�;�FZN�|�L�Մ�r�u仲FƦI�^�/L�X��� �O^�鑿�V�Hp�FD�B�Z<��F�:L���ߕd��I�|�%3�6MF|�PHe�q�����8�T�_I=Z�A$����j׫h���>q'o������UO�G��7��}�-P��ڨ���t���J+��S���ɸ��d��Mi�e��h8e1z>ƿM�JO�	�iX��{w���'߿кf?��/s��JW�: l|u�ˠJ<T1m�n�emO�V�e"E'���G�X��U�R���n���[x�ؙڬ1�W�`��c@��3K�r��gsȔhof�w�䰜CJ��uGFl'n@H�Ȩ�@�?������J�{Q��h�T}�g�r�@i'F8��v��Y���X�LH�����] �"x��E����g��K��2P�2w�QjYS��{4�?ɇO��<�V��vЋC�K2�+~�r3�N�%F]�Њb��a� ��m��B+E{��?£ J>X0�w��#����^�v��|�P��XlxV64EB    fa00    2b80���9�5�����ޔ�7Wb3Yf�@�^���:[���"�^ֱ�b��k���61 ����*a.�gPi��t٥�0��cM\@��l��cD�RA���6x�_�"�i�6�nŋSx���f�sY�v� �^�rK��hc���>��~���X>�6�T��Y�\�{t UI��0�ɂ�'�B�lSR�;R�É^Ӣ�:>\�	R�G�]�
X��J�'q;A}�_w�L8���4��w2O�ۿH�}�_^��D�W*ɾ�1��'��\Ě�X�Z����P���d4���=2`���.0�jA�h.�`Ʀ����pK�7�N�G.��rV������Ϻ�w�o˄��,�j��Y`�z�̷�&$`��q����Ӵ9��Ĳ�=�TU�W��1a�N�������L�W%RE��P�L�~7o��X�W����!c������q���v��geᣳ� ���C���sK�3�o�c�g�x������-�`~�\##�"��a�`ӭR��t�Q������e�E�������1)�+��]�g(X��tS�I>��et��H,�?��PI�.�|�P�W�,M�w���²�?�Yt8.���lf�hQ=~�L�LJ��c���)��K�%����Q}{�}꩜��4Zm ]����b�zS��@Xk��Qϔ�!k_�X��^��݀��r��S���ZQ̃F�A`��hYBG�$&�a<5�`�P�!�w��q/C�i��16�F�U"7wߥ�0<���%Ate��f����~8H��I�xB�d���˝f�p���Q`�e6���ʇ/щ��C���DVፊ�#��A�caY�K�Iӯ8�1E�g����f�j�.��No����#�[��7lb�B�Ě�R��O:�T�r����$���1�3�>��	Vx0Xw�G�̭��;ԞuwV6ʢ`YN4o��L�E� Ӟ<{`��~SV`�`�&E8l{F4�O藪"�E��"T�f�3f XA���W[0y�����P��倱������D��7�� q�U����׭ܦB_���MN�dYY &�-��3z���p�P�=۪X�������$K Ê���c�p��΄�����)���������Sܨ�U���ml��T.H�s~&r�y-���G���ǚde�:�ۣ�1�Mb�0X7��e4����==��m����&�Ѕ=��ŅÁ��y�u�o��J�t���\W$��x�D��.�1�\�M�b�E�d�l��k�%�~08�'�̡�%����3���COH��$G�̂@��ハb��&F��)įSP�N�ϗ���-U�fѴ��d��%�i�h��g?2����U�r���ȒG2b�LD�,�_�&�0գ�a�������a�V�0�0�,���w��T��QpӎѿLjS�e"�/B�QZ �'o�7�4x�t�mXN?���%N�-���ս�#�qIm�4�-O־X��(��k����%ƪNK���<O�X?QN��ɹ�ηQ�`tT4p�7I� ev2��Zy�sv����Kduл8�W���Pb�����+�1�[�W�z����>d���������c�������>T�	�+����	�� eg��e���0��g�Ӄ����&P|D�T�L����7�j��#�.'���.�wp����T��W9Q2�9�!�^A����v�_��g2d�� ׉����`���/n�rW�Iai�F���rlz�ds^�{�:F���+��>`HL(~ܪ�A�~!!�j�:Q%��5Tk팗��wĿ<�I�m {��-�(��sv�yrT�ݜ���u;�`��&�t��,���R�/�*��Z�'M�.�wD����a�U2�ޥ9tX�I:�oy��g��i��n4Sf8B�{�\o�uR���6#B�#�	�c����\D;> ��ho$���S�t�?|�H^V�.T˛�nr��.s(B(b��b�(�L�⋨�#�-�2��!M�;�5�Wj��V߸,%�߈�����Rg,�?��Db��k�6 5K����y�=�!t�9���s=�A�.$���W���o��;���QO�ބ�:�D��9~�����;�rw���"
�'�@��M��$�����:H긅�Ҕۚh!�f�7����X���Y�k��r�KW�RE�/L{�H�Ӵ ���$�%>B}\=\f����аsq@�B\U4z��w5���
H%ݽ����n@c;;�Af�z��Ar��nK��#�vy���d�h��/$vGC�*I4:����A������W:�y$圼���X�#'�q��#@�Xc��L�eJ͎p�'�Ϩ&p�[$�*���
>���d;�K���§-o�ޥk�Js��N�����e8�;,�)0n���m��a���g���=��k����_���_�8X�<i����K��@N9�ԦQ�tM
�F�\.�z�p�����C �4̎�݁��Lx�%|�N�	�&I��������	jr�s5��2�DK�x�Rb�%�N�9(��D��Oc��rj��X�Y7������e����$h�r�}v�	�#|�<gك�({� �N^��]�!�T�R�g�
�3(���\r����Yx12!�b*��duHq� ��v�S�����f�o,�h��Z�[�Z���L�!�(����!���?�>L�"
����,!¾OG��P9C�[�T�\��
Z�������l#T��&I�J>ZIm|F/nF���c���7�1$}��*�|�a]��{�@�B�����O[���l<{��u���=ɑ�/ĶR\��a�U͛ �AI5�( �F�k�L���6���Հ�T�^�J���j���~+��^G�o��l�:�"��Ms3��['�����@ ��"�l�+�2�����x��A��<��+�j	��n,�Ē%�9O� E7�#�:�1�J�h����a3�Y�^&�b���4;+����?	�U�M���hs�$.u��GU �<�z��x���$g���/jݭ����?Q��I�,�Y(��,�t�!���|&F�.���e�A�<^���*u�B�v��G��#jH�N��;Ym����)�8.3�P���+�

�y�!�%���~Yq>x�l29��x
���.s���3�����J��-Y�f��I�^��/��L��HU�?<˲��˄Jr�5�����/5��n�\�-�`�̚�{�EC�D�A���zZE�y��k.��1a�.0��I��Uܜ�GIb�e����=a��� u2��}9F{��������>b�Nӈ�LF(pqlu$�������G{����[��44;�V�rE�Q|zԌN�kB����f��@Yp�q�td��?�@�ȑͭ�
c��jEN�����������LP���0jUM�c��_l��ן��\/?$�+Jх��|Q�LG&4����ǣ�x��sW�s��L�9U���x�F��m���`L��a*�z<�<?f�����B����5~�/z�"���H�7�M�j��8���l�]I��U�MW�B�:7�)�]Fx�P4H��K�	�TZ9���`t��<��OTrS��koOVb{���-,���hF�bs\���y,OSN΋�$(�r3-Z�w��o�0��u�8��3���B��a����	����Á�>��)�dp}i��i��#�]�=X2Oׯ���.{DC֭ꋷ&�9���X���$���7�>)f#6P˻���d!1�杽�)��%w�]|fg͠"�զb�-Ɏ:�U(}�����$	�*e���R�d|�eǴ
���\��D�p���/��3g�5JgNI���qX;㶰��y(�Զ�O��֬����nc���Jl��Y(^�C��S�+	d��~�s��~S�1���/� �c�Έe65g�������cp��"f�5��r�`0��ȳUcM��r��'�­c������/0I<�s]�,U�f�J�ә��&)+"'=)W~Q+(�.���̾�"qT]�)�S�Z�7��j����}�V|�#��T�Ֆ���W蝭x�3�[�J��qF쳝.]]�9l0?��ʅ�K�g����� ���,KW��iHq��3�r���7_�KoC\F���Q�X$X�{�:D��M�^�!�A@��U�u�Y�)e�O۲u��t�!�m�켰V|�t}����4]C럗�Hͮ":�%|<�Q�ܛ�����	�F��]��'����g&1!d-E�[���@C[� j�W��w�,C2�&p��^+p�#xBf�o�f��BR�����:��gAy��
R*�;�@���6U(�Lz��(��3��'ޭ-�꣟f�s�/�qߖD�T�	#��ua_����~?J�*ux�Wb����,G+/?���[hT�jgj���~I�.��Isag�zv����]���>O��*�ԗ��z~��� _�������e9�S�m�|��pa�ʋ�)�JR]/��ڄ���:�'*�W��H�x�ݣ)����
�KlC�5KA�e1�Z�:Hw��36 9��0!*�M�/�姴w�䁈J�fl����խ��q�o*"��Ԗ&��m{5�9�D�PL�8#$O��/anI߯��xO�N�8�W!��.�3u��?�T��/�C]��}cz���W��<%G�1(Lx�r���Lbŷ��"��ތ��2VRT�վ��>�|L����u;D���z�0_
{��h�ƕd3��j�`n~ٵ!�>�f���c��A��Y�"��e_qMO��y3T������Ќ|�i��6���]J�㺔��x���5���!Uo�Wf&�.�U��9��C��R*��2z�]��P#�8�7J�a�N�!�C�8����_|l�X=��3"�q3���}���7	�'o�Qߒ;c��U�'xZa��c��>�^�_^��ѱl&/�%A��+��j�ڵC]��������^�uHB���O��2ބ'@QQM��(U����;��k��-�k7���Dz���r�q�TV�[|�8!w&�nߜ���3�m���-�,�SL�7���\[�I�<��q[��3(f�o��4Bd�,�2Fl	Z V�����'��<�O,���w%y*i���� /j`��(Xu��w#�~$51\�K��?��末��}��"��
$�B��<NXeW�� �/�v(���K�ejO�	ѿ,Ō"���c՜<ԊD��2�O2���0U��'��2����(��AL����(*� �i�������!|"��6�7z<��.����!(��-SOC�˸ȕ��Ǭ��ҿ����6}0!VH,ģ�%��?;+�dgp�}S���ct�!���'#��p4�=��� Y~�@����:���R��]��{��V�Nӆ[���>s�b�� Qg ���
�+�I;}��ļ��]^m�3��!��OF.m�kBi��>���X�[rH�w��@_�w�|��3� k�3�$��B?����آ��Dx�q�op&�K��{����� p]v���ƸJq�qZ9ל�����d��o�����<3u*�*++�6�p�Da�Ih" t�\;:0����/�|U��h_�By��wF�1�D������� b�i ���~����V����"
�$DVŞҰ��1;r��`��9����M��y~��i�W��
����h�g��D+����%��-c���x`�~(�U��ܑf���	<�!��3���)Nf]�]����D��銕n����48�,��Tԯ���tG��:4�1�	�K�|Q[��dJlhP��"��:�8��Ԙ� ��������@L>b;��F�n�>��9� �W�Γc�j��F����x\-A��\o�Wb�Ȇ��,�L�>c����g�܅��t/�SѣD��t(a쳨;7�G�!�T"I�Z�+��'��|�!h+�o�6G�9�ՙ���h�������j��e��c��lT`{�K�������gI
����k��%��7�<.�Ό�C9/��S��7�P$�	(��<`���m=�jc}�\�2/���?�dG��wO7��u������4�6��_��@��Ώ!�����t�~!�-H-�n��f
P`��M���\�	�2�:�����"��n��Q����FL_m���M����L�K�֪�������<�E�0��c#�RXy_Z����"�g�(��I�l�ڙ@!�޸�b�9!�'VeI�V������&����>�M���-U��X�\;��y�T^b�n!9v���y${��*��m<.�+x��x:�CQ����6t��r����k�����-����8�ݦ�w+��j*���Q)E%L_�]��TQC9��Kd���^��=O�: J�L����/u��"�k_T)UI[$	$-��`��Ϊ:;��)?�2{X�؋U� ������(p���q5ؙ��ff3a	|
��&����t�{=�\�f��{q��"Z���J'T�@�F�nB���0�H�n��b�(��~�����«iK��vKV�FR�������J��3�`��3Ϭ���JuGy��C�{�d�=��ڳ�V6�$��I�E����S%�����G��_F�d�:�u!�V�]�����u�(v�V��� cS����G��),�@����o*�x�G2�#�&���C|-�zw��B��$�dW�Q�����S��9A��<�j'������s�������Zd0~y�?d�R�$����҇����Ms�Jf�錷�T
��R�З����K�-N:ri�]�=�rM1ɫ�S=p�����b���(�0❈��>G�V,߬)�&Y�V�q#�RhY��.�����p���e���w��*)�@�l�꺷��g4&�\�G��H�B��|��A�=�<��R£Zł6�}`�o���vp���X��Sb7a)�#���B�Tj��M/�uM��@�!�i$��Elj�R�`�n;��^+.��{{����ڈϡ�e�ݓ�+D�\�jCz9@����Y�3�5�b#F��%|��Mb� p&Pl�l��6���M���"�Q����Ζ�H��ʞ� t04��h�O�"}�ݷ-ŝ(�QϯV	襈.�A�������^)@Fd�r�m���Nşz+[�r,{Re���D0s�Kwݒ*I�q:A�*��S��S�1G�L�0��wR,���OeNu��+��̞2���A�.:l���ƶ�N�Xw�Wc%]X�*_s���$ƺ���!Ef����L�涚��g2uę�(�����,�ceQ��+�1}�ռM�'��(#�BP5g�g��j'���&NF�[��W�bb0G�6Y��hn�����=����a�ۿ!x��6$���2��k�NH�����bv��oUU�6 ߭.�![�CDyx�ˤ�2,�?N(9�U'��}���
�J�Y�3�#<Ď�N	���#��,Vژ7���rF���[z
S�_��Jj=aBҟ߂1X�]�s:�G ��w_P')T�5����E}��įfd�HB���;Hz1];�*l�.��������˼����m������0;ݭ!��}V6��}��U��|!(��)Y��j�pQ��$�����{�t+��1���-�t	*r�
�[p��y���D;���M��ٞ��!|22%�q	h(����ɇ��UXd�Oꨙl��0B#v��b\�x����Y��Fjp��i�G�|��y�%�?̟�g�\W7���Ȩ�+�Ը�����%���[�,�`}L�xP��
;�:{�K���2�J;sÀ�b���IVl�@19���;�,� }�&׎�$?�tBL�a�EO�,���S ���jؔQ�e\��ѧ��<�,H��Lúh�z��J��i��I{@��!�)��
 �G����L�L
����^nȻH�n*v���(�C#��p�v����Q�zU/B:�vv��}|�O��`t�ߙM���C����e�X��\TI������U�	��r�u�c�F�<�v�nH�c;)ۮ�+��}	w&n�X�C������dm��H��c�����"y;-�>�Gmpq��N�����뤱�삕zAߠy�6^v��1������(����+�98h�+�m����n� x5}���WDJ�|Mow3T�2��7���h(��Q�l7�\��5�i����+�@��8[]p�gd��<v��K�c��
��[�� SF�_>����9����T�ѕQ��fW�aAH>C&�ZAņX9r�O��M�/���sf�9��j%�̢�雐��'�/��l���&�֌�&!-�ōǞ�W�Y���o?��h�th�w�~.��]y^�U��b���s��V�@����C�%�Ms�;�v�p��g|8NVu����]���!t9�R?��'�f z��Z
�/��{~N��=�!A�Q�Ѣ����ڧDmߊ&�[�����"�0O6"
�6�Cٛ�o���-5��� ��Cbp(t�J��Z@�[L��t�t��LX��Ӭ~8ߟ����q��)�(��͜�mM¸����#u͖���76"׏��x���	}*z��W�)�.u��s-2�]-/����S�����%_YD���%�rL�����$y��%�_@�X!k�V�;,l~`�����WAʾ�@�Y�ǠA},OF)�so�ݿ�EH��y'���E)���������I��,�I	b�pi�v������]> ����8�����A��L�yq�A)��!\��p����T���E�u��1�96U�E�I�-��[���<O��8������n��dY������O����Yp��R'�	��S�:9�^�j5V��i:���}�޳>1����9�������7x"�41�f� Vl���^~�T��K�&��"�|�ަ+j)9�4%��<d��w:�z��X�Ò�\�[|�a6r����N�`��}����!���d(��+���=%b�s���5����l8h"ޞ��1#�v>��wp/�k�f<,h��	.9�GV��t�E9�L5���&�e�"yiGv�7��fbw�	I���v3�e�%�Z�8��ϯ�kG ��?�X���|�1�/�dw�X,�u��8�+�����L�1�9��(U�	cLStbֶ��~-�ڥ��^�m���2�D�'�k"����s40��)\��_ t��ru.+_̚4L���ט3�b�E-}��!T}��
��&�6'�m ��S--����X�`�i�yD.=��72�&S�F#a�3��8�0�^q�}%l�J�lav9���5��<�:b�2�����f���[�S�U�{ݑt%���Ҿ5r�C���1(�z��w/"|��s�oO�N!�$��W�o����~�p���]�*?<���3�0Um�ͷ0���6c�
��굟S���2�E�@�C�X3�>���V��	���rgF!�9(x���a�(�X�@���]X�$�F�G�E�,?�����]3P�7h������|�^�%бpR��[R�uC�{��o�BԾ7Bϫ87gc,����V�N!��������{���Q1?�Ǧ�jzR�<��+6���ۈd���LŃ�ߖ݂�%�0O}�J'�lq����51$j挱�V����ٹb\�2�9u�0���qC���|�؋�q�a7'��v�� -�GEYu�Iϒґo-�hv���+���;���S���k'�]\O�E3s+�^�\ f��-0Ȝ�
g������2]�3��c�#���Ff,��Q��!}B��N*t^ո8Կr^�j6���ƽ�,59Vl���#� ��Q�wR�A�v�COm�qH�`ޫ_+��]'�"��2[	lCR��<��Eʓ�&��@��|�G�֐�ߖeu�Ҳ��y?n����FP�P^C��W�(��E8/��W:��z|z�(A��� x��''	��s�Z'���;LK��%[/󆆥!��
�g�fs޴�}
_��ÑFRV�GΒ�5����+���|<�t`��^����k��e��US������� k 
�.N�*���4o�C�ĘH/����  &|��K
��d�Eo8}�;�jM6�v���VauF�~��cmdC$�s����<�꧱���vN(��a��g�$� ���z��?�y��C��(��i�>�o(�Ё�o����PLnec4��?���*���?��2�q���ˎ&��(E��1��.z��_�h9���B �O�5�QPͥ���}h��uȇ!���͙9NH�7�u�� R����l�JS7Y�bEe�4y$E��1��Ã�|J3xF`?���^�6�E��og���ƽ8��*%J2Gt�q (f�M��.��ɾ���O�,U���*�>�$��M'&�/P�<DAEd��a,Л�����Q�B�_C.�b>�����1:��`���T��,v��Ǚ� %��?X�	�l�hu�܋�!+ت��Vl�aWqS�NL
�[��&�m�[e��3��dx�T�+x��Xj��֩�d65���Rߧ��lsk���zҢ� +e6�;Ͼ�q�Pr���(��bG,��<����s#��j4@-�O��b� o�S ������t� ��`���l��O��:T;�qܝ**�w�Ie��d�m���Q�>f���[�H��D7��v��~��nJ�D4��1Y���TQ9�]�6���R"�q`�`H8".����j�ŀ���_�C�ӁνF�����jYj���/�P�Ro���t������c;|C6�[�"j~��L��7H._A3a*�>�?O��z�T�qgg�F�� �'���z��������m��m�������Ɓ��7��N1��[YԊ	q��L�j��+B��:syB��@�c��}	ƭ��-�[�!G�^		�%�!��R"���K��ǻ�_�k>�Z�0Oq��э;n��S����*��S�� E�c@�DC�Æ�6uy�����_�����TJ4��H���袻%D��}�XlxV64EB    4ae1     d00�	`9'�%L���v����}�#���d�(7�Q��Y"܊�z���  oJ-",hP���M�*�`���w�e����ӹNb�V��j�D�:ۿ���6��j=��
�E��<UV'A�f�k��Y��<i*A	�	����P=�8m���!�ә��Ӌ@�w�D��3q��|��e�5�̦Jbx���c� ����1TIa�EU��ω�����EqEZOZ�ʷ�
��V��%R��	�C�K�ɵ^>��0��l��u��JՖ.�\2 �ל@�e�
���u�x��i�,����p Gz�90��$���/���}�Ё�}懥�[D@d�,!�/��{f�����!X�P���sfs��Qm�+~�2-���*���y���f�!z�9)ei�h�P��HS�,ڶk�`l]�9s���mۂ�~��@�d׮y}�\=D�
uK�b�r@�|6�!���*�2QX�dq�����[Kp�P� ���Ů��Ү�
�
�ę2T���s^%��$�0�_�_)��5��;fzu�sw��|'v��9.JK���c��K���4���Or���*��hA!�f7�R��ʂvM{"�0����"�����6Abͣ��H�����XB��͋VGs��%~�p�ٙ�x
�(�{ښb����D������Av���_��r�	4�ҋ��� +\8�6k˻���R�3q��Lw�F3��>pLC���%�<5^��$G�.n����!G��|�\�l���u4��MT�[>���Lj�a2$�Շ32"Xxth/�;�����K�F��9��$�"ܟ���X��cc8��k{0c!O���,�v��-t� ���G-�{�4`����zQW��?���%>��<�U���v�0fR{�LP>`aAI���*�7�}(n?(�oV�j'H�$Z�Y���]�P��ўS)�v���&��G��*�\$��[,}��Ԕ�j��x�\��~ќ9 ѯ�1t��N`�z���^9+��ֶD7��> �]��8���|�yʉ��S�����,���j��+�f~���4��°�9����$�n��ȉ�i���o�Q֣v����HrŃ^w��уA��}N0صW% x�.q
Ѡ?V	PZc,{�ͼ�����j�w�C��F�bNo30?x�;+�*7ڍ� ��(E��'Ϳ���o�������y��|4m���������;*o|Iؗ����M!��pČ�~LKni�so��j�]���DM���+6���|6L�g�~"}d:��ש��z&�E~��X?ys��@WV��ڳ�KL��J�UŐ�*�c�����G���7��/˾>�trKvLz�c�ǒ�y��_\	Y��P�J��Ӹ�#ɘ�3��|ݰ<�9���И~&F���4��J	Ի���&��Ο��[_L u�p�X�#�]���g��i~��:k����,�H7��)�W6(&��0�7��+,�Ym�D(��z� /���_�W���;0�U�M�ܳ~�wHM�e��k�#V�iL[�ٞ��`*W��l�0z7/SAcydIL�0��RP�4��LGLw2b�m��D�*T�\;U�gpݙm�3�Rt�X�}*¦|D۟V��Q1:��1g,������D���!+÷�Z�b�F���/�����%�A3��î��lC�մVV�b8�6�(����,�d���Ne���@��\�o�>��/�d�ogjMy������Ĭ �}�)0�����L�;-h��g�����z_BhO1�F/4�U�@����<��f��T���f$�&�/|χ�OLg�XL�hޮ,F�4���V_a�S���}"�i"wpG����FR�֭��c��s0�����z��S��e�m����<�45����`Sk�Y�.�.��03��s�V�ӆ+Lu�Jϳ�!�l Ҵ�����Т��D�	S��]�y	Y���T#�cң�z���\�ʡ����r��Q�����:�?���+Y�|�Y���+:?�9q}3���m*.N�I��S	eNpPɆ���,�d��(�߫�xy	�u�;ۍ��P���}B�t���.���"QIS�;*��*k�UO#�u�h*.��qQLB��Pf�/<�D����7���1G�u����		��Ҧov�±f א��E\p@��?\��������rGnÛ�H��[� 纍���n�U�����%���='F1N�mlmЭ��Զ�K�TA}Wv.W(D-�͘��] �-�mڳ)���u�D����� ���r���V�9ބ�p�X���=G�V�z�֚ꉯ2Օ���c����V�wC�gzyq�9r���R���z��E?�I,t��.f]	�����!���N���t�ZC�Mv�I#:.g4�(�E��͜��F,���W<U.1���h�?���;�P�|+������+|�������G��.M&l������h��Q_Z�)��]"H�u����3�5�p.U�׉����9�祄�DW�7��<�Z5�q Ę�d�e��.�hHb��PL~�D�a��nS�|��>�:��mC��@��� �8%��A�{(�O�K���3�~}��ϼF����<Y5@l!ӕ�B��Y�TDY��T1�?0�����$^8P�®�o	�0|*@K�Č�'�I���rL�a_���J3����!�nר�b&��2��jGQ�y�.�k��(Mw �B)��܂q˻��kXs��dbK���!��-II:Z��d���Y�Z�t�Sثa��6ډz�U[�d�S�85F�:�����9;�D-P���p�(.��W�R���e�B{��Vm���,R1���
�gG����
�J����p��h����Ͷ�ž�����J)7
p���}W2/�1��z��i�[�����i��q,6���ɝ_�-��$s ̖���qFS���툼O����(�.�ٿ5ڞp�k�A���K����F�qN��S��t7h%@�h<]��kRӒ�:g}�3�	��<��z|>�B�]*%��J�̌�P�_4�f�5����b�d�Y}e���K�� ͗_4{�3y�E`6�D��O���=��q��mv� �)��&�e���׾���� LU�K)�9�̃�:lMS����M��@��y 1�)�xA�_j*e�@��SV'o�Z�V��ɷ�6c�3ƣ��B&�ު����t��]�ɺ�1WN�\�ax��9�?҉����m�sn�����'X+�6��'��5��5oEX�H�^j+�Bڀ~��r��qD