XlxV64EB    23a1     b30��l�%g�������?�Kr���OUwg{#1nN,n��a���U���
Zh����]����R��n�����>�/?�-7����8Q�t�V��(-���rؚQu �b-#vG.C)p@p�tT�AL��e�#+����x��l���"���o���{����MS��Jj�%���f�4 n=�ȓ�E�s�����ݥ��&384�'t�����2�@ȫ����\���K�_����6��n��-�a�?�t�0IU���a	�uH#�N���-���D
;�u��Mº��H�)�Ş]�����T�k�GH&�қVܼ&��é���s����}�^�2��k���?-�>����N�T�g��xm�����ڀ�I/0JS�c/{F�BO���ߩG��i����B�`7�/�m�ly�O�հ"����i�&J1��!���u�|l0+H��e �S�pf��=c����0�~8���a�]W���3�0G >s��C�<�6�zo{\�X7���c�OIP~O��]�!��{��^,�h(K�[��	�e�W&pSItQ����ͭ4���Ц.�
�ˇ�J㮭2'op& ������ï�.窛>�[�i��Fy�y���pf�&��#	3iD�APB`JG���	'��?}4��G8�����7�-��T�~���-Ѡf&����;i���׻��J�a���(J5��D�z���"z�frk��f�"->�
�uU���KІjM����W��_Ijc��ǹB��yGAږ�u��	Y��6��dP��n���P(M���hm*\�S����49�S|׭��L[�q�j+�����m@�i�x���.�"E�e�~3�'�瞰i�>c�r��A�n�h'� qT)
]�N"�[iR�k�ݏ�*�W�����J;̩��KY;�W����!$���Ao�.�&�������"��I���g���=��<�Iq�UE�[Q;3��tʍu�A&c��CT��7װi�f7����E r��ѣ��6��G�䤘ϫ(�S�(1 �~�����p��d�|��z~i���
����L�>����*Q˻����h;�z�'��s�#Pk�,����2���"W)�pC-�Y�	�0�[|�M{�����"�C/���7���M�	�����b־ �m�H��gj1�5R����f�8,ڏ��)���Y�ӑ�K)��b���E+�{'�2kͬ�$�^����Q=���TG%�Ҍ����9E�gT�5T�
h�.9�����m���t2{{P���ĥtQ�ג7����e�Dx\��;8�4��NHw־+��7���Y�����1�;Dd<���<�,E���K��]7��
�>q��IKY����U���ǿD?ݗ/t�E�<��*�+�%H���_m"�Y�AW�ˮޝ���2u�w�o�����3�(6���G=�� �$% �Y������s���:��ܫ*�fC]'I.�Q��v�l�)��,M�����D�]r��ڇ}!���61���e�}`g�К�j���"+�K5�f�����8�.s'
������nlD���k�}�� �1�ʺq�Xy�p� j�G�C�g1'e��Nef��)�(���l�.�NwąM5��XQ6p���aq�xoa���r�q���$�dJ2�c.���I0[[��w�\k��f7��u��d�u�gΐH�����K�Wf��l�Wp	"ɜ�[M����~]��h\�y2癢��fȶ9�m�9Y�uK��{��.{N�=���������pIaw���fV!AO�ꈺ;���j��N�L|�w)�	�m��C�d3����BDfU7X������Xj؊�=���T9h�,���=KklHx���(+WW����{i�@�ln���0�U�&�����{yt}�>��!;�	�~=�D��P�
%yNP���	x�ju�(�� ��/_?	m�5�k�W�v�*�Ape-N�$�TL�*��Z�d�v���WV���_�_?�o!AR[����"�k�z�(H�;@���t��+�r#Bփ���qo�a�33{O	џ���N�n��<�2#�u|{���=LCm��(�,�D�zz?��L����������S���]������V��6��s��/���d���V��Kq}8�$�7�+�u�)4���j[,�� �>@$�=#-�A�YB���%�T�Z���e�=?A�U.�c+pfɴL�#01m� 9�l���C�Y�fm�?-����u�l����GZ�&��^V���FQ*k���3+3F�X��-�� !�D�؀��uo9����H7fx^��YgL2.Dy"�Dww��)��R������YТʇ�'�u�$Ձ���
5����cZ!^R��Nyl����?o٪�lc�,;�$lE�Nk\�e�)f�z��pj&:^��Md�^6�+�A�9�gw�5��H��9�r��er} N�r�쇭�{��~���K9����S����@z��O����0뗇�om ���rEp��G m�jx��mjlܼ;�'3餀t�i����!�^���i"��<qn���3�ݤ�|l��9���q?P߉�h���o����������	���+h	[(Ga��.?1�fYO���Ev�\��?�X�Z�Y189�b�X,��Z!�|5�1N����[�{_+��v�{�����;{@$[�2�*�on�7ߙ, �&��Vh��0�"�w34
�*H�=3��3�r��Wx`�����̍�tvA�	PV~U8^L��LQ�X��$������=���dO�d �9�3h�Uf�|�o��L����b���^��2��
�q��aA�G D_@�9v\�e�23�0�IGZo�%��M��x��Ia��