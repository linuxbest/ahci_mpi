XlxV64EB    24b0     c60UJ�?_��X�Գg&J<zܽ-������Ea0��g ��j�@ۉ�D8mes3���(Q,�o�_Rv��Z���l.b�VJy�]��h�R��D���?��YwX[�姘겇y)e����y��|߇9��:�n���V;S�ש����.��9Q|@[�-���rX�f�ڀФ�� =��G*�9k+\�4��N�>6�ϛ��@Gѥ��L�֒���<�D �;O�<�o�4�oʹH&�c���?�pA]5]"���h�%Zjouy{��*
�T��qx6eJlI��z���V�&�pR��d@������56EtK��\G�V ��(�_�xO����g}���4Y8��j��\C��T�x^ ��6 ���j륊b�X�p���p2^��U�8Ƚ%�H����{;~�A��qd�d���5L�x[Zِǵ���3VB�"#+��wF���ET��
�d���J�|a�u[��CE�C
_���^e
#UI-���$)5���~5�.1C| ���J�>��V\�o�*{�%Rg��?X�%ߌ�&�ʼ��D��az�[u];�����D\�i�� �<:�Qp�CBwM�w�
}�J�Mh��ej��*��x���ˮhS�:�#6�����G��C�Iʹ���R���ҩ��7Id#���޷�S���)O���G��X��ҰY�u׆�&_��;ĘaN�z�3͸Zo���P�#H���쌣u�������b�k�K�?�C(眢�I�{.�On� N��Ƞ�D�^��-yҔ*��H�&�4J�K��cT}�P�u����˨_�߭� _�*s>с\+�z�^��^��0؀$��������/<=�
�z�[��$}��!I�~m��	?~�G��.NΉ0���V�,���-Ik�+��Oʊ��Q�H�%.)�w$���q��ݎ���4�� j-f�>$#�&r�lԯ8�S�I�\*o������ l"�F[�1�J���mY�""�1C�X_����z(�G��f��}S����ʿX�V�Fz)0 Tn���k��K����6JmJKs�V��ȍ"������U=�	���8J���}�@�r�S���qT���Y"Y��
c�K/��J�iO,:|�h��a��w���A�S�[P�:�~j\��?'2�	M�'�%sڮ^Kt>d�n��4z结��ÿD��w�e�X8�Jz��}�"�,��Z�Q{��ZG�MdV���1�ͣ"Rb�9.����&��
3V��d��Ǜ_��KG��7��n�QU,��}��c���Z���!�B�SGg���{�S�U����ʺw6�1�}ZϜ�^��Q	��ns�#��Չg,�)�Gt���M�֊�r�p�'./�oUk���&`��s>>:�K�PL��ީ��nTvT�ͳ&����{TFGW� ��1�^k���[��_�L󣆻~���y�[S�:�\����\�s���w���e��������|4�ُ-�W:S�1^tt��wJ�凝�<(_��Ȳ��4����9s���}?PAm`���uD�βg�e�`n�<ӄ��Cu�����x�������)�u��vc6�s0�����*j[mJ(W��Պ6Z�r��	�v�����?�w��Z�У$[b����ǁ�AsR���Ч��S�OH/�%k���v�L���N�f���1Pz��n������.�7�cn����ܐn���mOO�q����WʂU!#�/tqZ8&�"޻�- �S蝂܍���Q[n�-"����蔕*s�MTϘ����?����=r��M��B��|�E|��-�no�E��a%����2����r����<�T��ȡ���a�h���+`ė4�R˽pX�;�*��Z�0ԗ:��}֗��rcg�\��y�z�`��T+���]��j��sr�V��~�9[�1���ҙ~-����PN��q�T�e��c	���q��UIqk�FΎ��5���b)�+�EjO�r��mR��E�I y�ej�\���bg�-�������hô}40)���G}���1��;�����	����/#�s�;�Y�yF�L����F��	���)��Y`�!������sY�U�,z��Q�� �B�D�2��� ����PA�J�,����o[#���Õ"�,����.enO|�x�O����{ԯ_X��������:����t������S2�udɶ�諀BFO�3IʫoM�d|��a<�:`�� �FQ�w���>(�YmEG�Q}Vlm���湱���J&%��o���1x��x�vt4�w�`�IZ| ��`Ȓ>��yvq6!��{]u����E���]�6��1	h��gh��\�6,����þ� �,�3sr��Mq9�n$R`��t�CS�W"~5	��\B)�����XK���䋯顗�[8a+R"��t�&$~iO��uъ�7�yt>ë�����9��9v(���5�-� S�y��m��R�{O��Fgc7��a���)��r�_�|g�|��v�ծ��-�J����Y��q��,�4W�%��6@��L2�<�}�6#���%�]l_f�������f4�h���|�)���ك]�c�c4��8\	�٭\����8҆o>Zq��
�����&�[�j�z-ۇ��%W�<zT�����절��q��܉nmc�����ܭ�ТV��J�� 7�M�w�xn�s�/|�Sm��z"Y�҄�È*{��-��j@��h��D?����I����|ښ�G&�q�T��_�.�J!���'�\t贙����>AQjϖ��i��1���9KQ��q_��0D̩h!��|�*A\�C1L��ܹ/��+;d3v��$^�v:��T$�@)�M|�#/h<+�eB�6��X�u��%�>[�گ���n�$�{�|������jK�*��b�S��'�L�RD���<��Q�}�.������Z�}<پ�d��-�n��l ���Ήc�_�k�ح���8�JO/�Eb���J�	4�����&o>5hV�n�y���Y�@H:�k����Q#��w�ek��3���8�� ��C�˵v��bb��WY������>��yA5{N{QC�:ݷ)JF"M�J����$"��!�-6Uqg�V��MT(&H�