XlxV64EB    fa00    2f80��L�V�=�H���b	1 W`n�(�.�)�[##,��R�����?Ad�Q�C���� ��_ێ��	�q�s����"�g��@�N�r��*̓m�e�D9:x���l�=�Ò��:�R"_oNA%���"�'W��ND�0���!�LB!������u��ƺ�1��ɁՔKv�Ǡ�O:r��z��Vv�$���={���ˡөm�,�-��L׽��_(�0�Y̝~���|T�"T�������T���<�pt��ML�jX��I�N(����a���Mx�t��� #��Q�/1DVm���l3P�*,�or�I0�G�0��ϗc������&��Y̱����6�H��������#����]�YN%�)G�A��qj���(�^M=���9x�ʯ��L*�<������*���!�bx����xg@ؖY�|�d�0I��+Lɜ�G��Ij��fpR+���Eh���9��]���;��>��U9!�T&��⁁Ǵ�:�_̏�drګ�Se��(	��f�h33�����ɽb!�Z$t����f���t�����*�*��)\�0��ƛd%G0�����"����kޟn��h���Y�Xܵxg�[��1��O������y��\+9�{�N[2�����6:�_�m�~�D�������k���tATe=���|�Pb)�pЅW�vh��^x�^ح�x�A��������l���[�)����w�4� E�cj�y���tS�퓟������[���yZ%��bL�]�{�?$p�Jd��p�#��B�p�Gh�Z�q��#�S��
{$Kq/��d��#������^�Hxh�4Hŗs�~z��c�`�z���ܓ� W��-�@�Mnv���3�~�E���7���Ct�.d�5�`A�ی:�ͯ��E�s�MK���g��V���I��+̻��e�T*�D9��P��'x`�	W\m��FcR��ʢ�[Zw�a�o?V(	
�Si��w�VQ��c���I�t��BÁI�����R4Jl�'�yZڑ�{A�P���UR-��п�@� #��p��|yA���5}m�f��	Nu�������P\���+rSi��/c��sMۇ;e[WD)����ak�lL+���@ ��,7.�Ip]�݂n�V�E��� *zl��N�%�!����؃�^��UL�B>�t����������ǯ��A��>����P�"��g�<�#@��ҜQ���)<W�>�߶� ��
]��/�w}���l0i{�D��jH�7c9SW��O+�bِ^��S(Vz�Y�⏌ൃ$���SجW�6e\����s;���d�c/}T����O�Y44�v�m+����g�ƒ��:�A�����O�-nOژ�3>�Ҍۦ��1,_���y�px��g������C�%@�F����L��k��	��Dڬ�Ŗ��d�rʵ��X��`W����e���:���}[/�R�e�mN�J3"���v�S#b��ZIzM�0�X4��ؓ�J���󡡠د����|��`��� lЪj�PdB�J|�	��l�o�`������Hi�t���(��E��<��p�LE�#<<���V�� *���W�@#UhH\�������:4P^d�j�6v�B3�=�NV��0&I>�����։���*/��!\�%ݍ`b#�52�5�d�\藞���┧���@���ҋj�v�ۘ���A�/��Okr|��E?�6*������p��DO�48�!^Qyߠ�B��f춛�c:7`~	DG��9�̿}OZ �{BJu�ɖS�HV�d���V!��T�ɇ��V��m3̽� ����<�R�.��#y��g�dq�hr;Y�b����f#m.�Y�����S�q���Uqؿb�� s�?{C{�yz�x�e�ksx��u/���;az�VhקT�c����u�X[�9aYuS���d�ou�T�dʆ^SL��Y��������1�L,w��_Ws�4� ����$�>Z
t�$�o}�;�������g�TʇxwE zb6��!�qJ<�,�'|i��7���>��D�]��O~�̩�VGρ��u�C.߹:|���"Q��Ej;T�o
t�qL!�L�雪��tI��5thE�!
��3[�ӑ�Q�zf���.o�c�qe��	�HDaM����I���_J�y�b�'C y��Q��p���5��n��Y�?��4����"Cbq`���Q�
�j{�I��aR�Q�Z�p	��̩hw��wb�H��f�z�#�Z��Z����R!����zI�wϦ�c��R�s�#����Cѽ���<WA�W����%��L��Cg�B��lfx����I拂7�;�e�t�e��3����^1��$ޱu1�y�F)K��nx�x&`�ޕBo'#sC�V���}"x�e����ij���Hz:H׼0�uW8�P'��ȐRf�
eX��LT�^[vsa�#��ٽ�����71(���kk�
e�p��9�2����)�-�R�R��h��o����nұo���o��K�%�ϑK�Z)�l�BՀ�K����t����HB�h��d£G��mѭTs�W~����z>�2S�x1�i���C_�0{l�_?uͫ��Q��$�PZD�1ݶ��,üJ��m���ƭS�d��J��kƇ�9Q�
�����Q�+��T]����c�C8����vɆ`�٧�>��)$o�V���q^�8�(���Wz<�&��a�U��K�i]���8��Ê�O�X��v-7 ��*����3`t����E��͝[��fA���J7��Ûj�s{!ŋtB�E���_�j T	�q�NjޒOI���-7��ݟ��l��_^*�;���ۄ��Q�,�]�6�C�|�������Vn��o`H��j{��ֻ��:<�k�]ˁ�BQ�����o�L�Ol��<����S�A#_�P�p�i�p�-���S��_aI�a����������0���7�T�����M1�$����!%���Z�~/�,��vjv�'�鄱)� �>����+�k*RN�#�E��=QtF{a#�����S���^����Z�Y��*Hy^����%�2B%�FIwzc��V��1n&��`�υK�U f�M {������?�+O����\J%9*֡!���R�PS��Bu��U�1�>��@4�n���:w��(��Ů_��	5菍���bt�8^�P&���9h��ʇe�_�����a��.��^�����s7�(W��As;�����q�c��q1�Kj�P��O���G�=���C����YP'`3�	�E�D�@�,�v���M:�I�X��i���-�/A��Q�'�1`����5s��iH<]kv�ԳC댩�(>?�*V��j[�G�sݚ�򇲢�
M�}��h��U�F%�78mm�[��1�B�>��m������"����N�'�X���!����YQv���y,4�*' ��]�L��R��<*4�L/���ӽ����ϵ��(��Y��9���öQ%S�l���}�����&ͷ�Z��Ω<����-2�(*�ui���O|>�Pȥc�#H���\h&��:Uۭր���]��7���B�����w�V�A�YV�S/�p`��Ax��S(�d)R@s��D]�opᝍn}�m����V0t��	�FC�S	�ٗɒ|	�L���^�����=+�O<�~wgfV�]��v�RM�j{, %��{�A��v���"�CI���~�q6��J����FlvI$k�`5ȡ�Ɔ$`�m�*uc�׺B��m����#�5f�j;ON�kUS$:��S�X��(ч���{�X�1K�;5P�sĚ1�WX�ڂ�h���c���/K�*UR+E�FX��x�b��Ԯ��罙,��#�^���/��Le��YJc|졛
b��~[���� ���i�'}��W?�$m�2�N2�08� 2V���0���γ���������{�&G��qxγ�9Fz���+:����AE.��֬��F�Lކ$4vPev��04<��US!�@��ҡ rl�J"�1>D鮫M���YU6��IS�����<� %&��80��e��{Ͻ������[�����	� \�M�<�p�m�q��*x,�r<�����{��#���/��RH�{ߓ�Z���"�1�~�ҷ�	$I�"�����}ӻ�K� �����l7�� �K��D$��ELj���x�s+����4%���Fi���(������׃��(\�{��)�č
�����2�t=!�B"�,�K��?�+����(ʦj���M��=l��L>8��ha�2�,C�����gA�ǝ�l�}f�(�N ���1��<Ԛ!�~�%�G�_���9Җ��Z]�h`GbE�u��kX*[)S��-�7� ��$_�/�����?J��h5b��l��j��A�x'�7X�6��Dl7�n�����j��"<nx�kdئ�E'���ZvO��	�Vl8P��h�m �T�5���}K�uįt�	*ڼ�ST�j��I �w�f��1v�]�b������G��	��4S9J{%%z(i8��S�?�SZ����NE�e+�ƔrβJ)��h�
Qa$ؗu��t�*�����.���D���,n=������-�G�����p=�|7���@86��ѐ\��������Xוd��������W��Y�B�Ȉ<	}��א��3�	9���B�fG�. �C�.�?���V�{�e���&1�.�F�d���x�HcP)~hW������tW�Ms��;e������=�.��&i���.���a�V��_�wdkX�I �S;�����O���E
"��Dl���hu�:2�J�����y8���%&:Z;l]�f�f-J��Y�-#4(b���Z ���n.�H` &m�\'�ߍ�7z1u��Vxc�%&�S����(�����)�>�;�c��g#Z��Z֠N)ђ^\��G��tN�� �m��X���c]e��9?z-�b��ߜ<���70�W\k�8��	�g�τ���H�ד"{9ւ�DL:P�nR�l���\�v�m������XJ+�ZM=&�Z@&}Cr�I;KwrQ��K �0m�YQQ�2��?�e���P&1V��u��!�y��%��:��F�WC�߁EΖY���vMmJ���XI_�ߎr�!ˍ��@.c;� ���z92#�$�[H���C`"�)���L[O�nm��i�?�!�T�*��R�9�{����x� �˸6�?�7V�`���k�T�}/g��8[j�?,Lڶ�����ܼ�tuq}�0�_ψ�'£����-_�KM~bϔ��4�BQS����E�]k>O|�v�ډ��σ��T�ǌ�����}�~IF���kdM/`߿El�E��1�dCU��T�]��2`���k^�xwf��L��K����>�*�j�Q�PkGR�n,)���5&�(��]oΑ��D�p�߻����^
gAq�|`��$)A��]���"J�U������2^��Ym�W��;$���ɬU(Z��tV��R�To�8�?�CB���<�Y�2���
Մ�Iq�{��-�&h�tq�[<\^��+�����L�L���İ�K�ɓ`P�KqW&�c� �'p�ٟ���J^oLm6Z3�4�"@ZZI��]P2��Z��18!O���s�����n���w�t����G�"�n9q�B��N�Li$���*Ư�4�/,��	��[�f���i�ܧ�3%�E>�ݯ-I����Z�q���
q๺iSԽ�f�m�y> ���d����$� ܡO�����W^�g��GA�8n��4ZdPM�'�w�v	�|��yL�d��}�<zy�
��+}Y��ޕ�����aU&>J����hQ&`<μ��A��b�aPFֱ����
i�4��P����lE���&�@�O��Wa��&�nbM���}͗l�6m���"!���c����Ck\�ݸy=?�d��dZq���,�W�	�As �Ss�����ns�D�H�0�C���`�d8<�iS�}�
��K8�N�g~x�UCL����W$Ϊ
�tF1%�B�����<,2���n�j�����B�#X�nT狊<4��s���xc�{l����#]��ۣ9�LbPE쾈Vo	6h	6I��d�Dt�Zu��ٳ�{͘�j��%�h���˝&�N�l�Jp�k�RA.H��M��&�5H�5��,����B�i�3ɻ Jg�q��S�M�0����E�,���c�	�a���mM�}���C�<j*�ۆ�"�*Ȉ��m	�1̃�KXRש�p�I��Q�ϴq-x&�ŕ�s��V���B���z��1<I���WƁ�W��W�F�O��g��h�0F����nMa�a8G�
Un��(����=�5ټ���٢(�17j�t[�-���?m�kc���a�$�5 ������YamxK��n��@�2f�G��@�+��F�W50YU_/:08��zߐ��8�x���h09��	��z����*�ۡiL�#�Z�
������_VM|g1LjaTpՠ�g23�<��������K�&��;��� y�0XϽ�zV���@޻��%��D�N�� Ҵ���kΨM�_���Uz�?Z؀_`�f�`����s����>�0��$� �u�|����2%�8M���*�"��9��VB����?��3^�_�XĚ�g)S��z}��kd�i�)��e�"�����f���sQ쵧�Kc�g�ݒ�V��5�lQ{�ޣvyJ��E���ڲ���5}��o�\�o�xg�ǡ#`�����x��m
/�?��	�%'|�Č�6�R�����h߶�� ���s@���D�D5ået)�o��\8Bc������C�p^�Q���b�^z�R��o�i�q�,-!Oe�S���D�$����_�h�֖���z�$���Cf��ۘF�2�9!�V�4c8�zfmdZ�j���&s�?>Z邯@�Os�����e���W��p�ˇd�Г��4'�1���̹x[ൔh��Z��8df�+s3ӄs�!X�{
�+p���R���e[M�� ća�Լ��@����Y���ڲ5�_�����	B����SK4�"����A��Y`��{��ssQ�5��G:5��;���.��[E`b�p�g�����dC~׌�e����{�>ۭ6H��R�:%��8���(l&����g��6;M�F����d�ox%x/
0I�D��-�' �N��d�H=R��n��V��\���y=�z���Tq�tn\.�J8���M	��ۤ�������u:��'�_�3n���:&�Μ��3����y�;#ww�Z	�w�3-"�,삝@N�wx�`(�N"|)�xE�G;ŅY�F�~ė��7C�����]�H�)x]���G����2�Og�F#��a����K@�]YLe���!���(�p�B��v�����7}T�J;����u�Tq�Ҵq�Ӭ��o�� >��%쑩X��!N"�+��j�$�����&�lEv5� ���dE�L��RN�q0���hG���㥸��b�H��1����M�`� ||����4���P~�ٳz�X{d�����9 �v/����Y�h���h��'�-HVӺ�P�z�^�I�TM?p GqŘq+ύ�F~W�+}����i��W7�U���/�ø��$�,�©5v~�UX�voqǖ�d]���c�d�L`��K�Ss�}Ya됁�@��s`��+Ԥ��u�Bc�~�����ZwT/4(_�1=\��o����=®�K!���<�(8Yv�S��'<����҆w��FÔ�"�P>�7Q��)%��4���gIR�٩aL>R���5�@��i��:���)��)���6���v	/O���StZچg�����dh�Ȧ�%#�<.{e�ZG����R��5J�H�)�{�P���q]"G�kzfO��]���R�d=M����4�)��/�4�T�a�x���E�ѐ�r�Pj�wA�s�X���h�j_�P���^�$A��-���\:����le��	����ۋ�4��z�t�>�N��(�/r�5p��t~���uؖ���~�4��_M^���I���{��M���LEh�q�6��a���Z�A��)��1H@D)1S�����]�Q�W%Cm{ʉ���A)z�f5�8g#���@�������x�һvEc	���ϝ�8`c��<ɥ���t�BgX�hq#���$��IR%�
��T��Jd�ջ"~�}�He�n� M��#�ۄt6jh�U�TI�J��͕FޚY>�.���S�d�Y��Z��W�N�˄!�^6Ɨ�#�$ۭ��B�(x��(6����r�nx�?�̬����2mA�����򸋅++����- �fu��L"��?�����4.�$:�ٯn։�Lb��Y�g!7�[�"�������%��qg9�U�0�}h�Q���#r��t&�$nAL:�:����~@`i��"��t=�����L�$��E�z�TE!��ףscz�vj��R��G�jF��}lso_���g��#�g3�����ү�Si�u%�8��R�W��?�ֻ��(�`���2�P�.���1������B��=8&;�:���K}
̷c犮�'�u�����O-vMc;�s�Or�6�D��;JW~��+�/�.�ʃ~A}��ӝ:��r~VÁ�hf�H��xj7�����.����;-6��.e��D�Z��['pw�9�����ɳG1�� p{�M���98����u!H	�>~L�'�qyj]��|Ð�G�C��UhJ/ĜI�C44��f�r�NzŸ�f���h��tC�k�+��b?p�ܦq�I
�O�;��Iu���ϚD���X�Z|l5P�����j�T�����1�:�G�sI��R_��d���mw5�3�;��i aNq�}����7[��?�P��g��ꈌ�Q%�<�Do V4`��x��).����Cqzt��Y%�h���h_�	���4�3�QE�>��VµD�
�|�`'��O���t�y|A� �pr�G;�l��A�"� 2b������ߞ\���F��A�V�^�k~?��o.�[)� �IjPA��sS��dОQs6@O�C80���Rh���>�X��w7pf<�J����l��h��VXe�� ���<��d6�i� ��V�{���b��V1=������ZO}x��X�oʑ~�2@�����oT�G�v�L��n�V7�Q��F�G��h�5�*����(?�QrA�٤He�$�
{����T\�䈳��3�i�V�W��'��n��h*S?����T�`6qK��ȌN'*J8���&�ف�X�ŧ�f�D-���8���_q�Um
>����xSa � JT'� �q��-���C����pV�"4.J�+O�D�Wq�K�֗�M6��A���S�W#��O�h�)� 4�Qpn�C��Y�'LU���h�Yq����R�b�-D[�Ld~L���Oy��j�]6�w�F$��$3
��+��Cs�+��V���K0Iڱka�t���<���yM�ǡ��?��gg�l{�\���
xu%�6� ��~��6�C\$_�E��B�<�<�˭��6&Xb���S��6֟�-�(+��&,b��g����%��(�>nlAU&�'rW�xiA,S�j$��Cm1�v���E���`���ρ!�^iɥX��Xty�1��z_��ٯ���'Fq=�v�3�g-e���� D}L����Z�����j��נ+����ټ��b��k��p*ԤS��>ť�����Moj8�ʹ�QW��u�&O�S��h�I�����߻L�D��^6!e�Pfк���)+pk�m��f�{DsiN�T�)�{Q�#m*3��=<�Yj(���c'�,��]�*����'w�݌�r�^o� @ןF���5��Ņ�l4����9�Uw�#��is��՜-C\�n�������_]d���6'��²I
hI��~�����N|��^�G��s�
}c�~e�K�qX��챬/!��P$6�躋�_9�2�g�� �������a���[D]<�|��j�ߎ�8P,�}a���[ ��a��cg	�
��<VZs�ւE����'���ڜպ
 �0��u��۵�	>侑��f -���̘��Gˇ���c�b�Rb��.+�S��4�3��;b���T#�,�|��4�0�^(�-&�4e-�iϻ,�T\^H�Rl�n-�@��7k���|[���.A�YD�غ-���ܗ�s�yv%G��#01L��M�r������ߠr���?�d����g2��V��;��U���.-�9��UnC4�6��k���s�Ӻ��ϾԒ	�ct�b����D%��ѵ;�lo�w�KC7��>c�N2��}4���E�0�s;:��� p��7��8,pG3-l�_F�pR���ϝ4�3�%�ޭ��V��~+	��U�9 -s�dm���R�|�aJغ:�^����[��E3����.E{����+K��U�B�����0�b���dΒmɩc�IsM[9ud���n���X_C�p]�bm�D�9���m�LR2nڼo9�W.���f+8�O�b���YY�z���4�%E�}c��6bSm�
̑�"�a��cr�Ki��Us�oJl�C����O'��uңvD��ǝ��Ӂ��v�4�q �����|�J�e'=�$x�)���qw�B1�R�ɴ��,BE�"��N�Yٮ>�vvvK�-zƲ\����1�t/�2��I��{B �Y�q�۝#�p�.��S��I�O�µ���*�g3�|����ܨ��`���eu�}/*[�7�^ٰ���xT嶡�G5��T��)��=�٣e�TL�`�#^�}� �qb���-�_�kۗ�p�%G���*���y�B�7_1�b���-enc�X��mx��|����-~>����?&Wq�a�%a�W��?3�E��iu�G�-��A��������MX��_�XG�#0��p�u�߭�������#�+-$e��Y9�Q��:��W!!<C@�Jf��4?�N����{����O�3l�3�ݺ��E�,�Z>�WֻP�n&�H�kBou����!�n�R��T첐�P�!�
/�ò�� ��Q鯬���~����5�ކ߃���>ӎ3���c}���j�.��k;((��P9m�i�b���	��2bN�b?��W?�p�Q���}�)�C�G����a���e��s�@�9��C��G�]���m���,30ΘE�Fv�7sU@���O
_����q�`��ө�>�H�aE:�˹p�X����?`��D��<����K'|
q@�jh�w?�Q��a�����C"\�@�">��Fv2�+��{��� :zka�%�D��"R1;�ejNH̆S��#�/�D�N
������.A���bOa�^p/�)�˯�;��S���DDZP�7q�Y�'�GN.!̉��l/93�wd�Ҍ�?��ܣa�_pY�wZ,�KeI_�0�܅D�[�Q�ĝpkMyE�)�O�%I_�Wݚ=L���h�7(�Q7̓+Ћ�E���,�WO�%��}�q+"��k�bJj"ڿVE�a^��K,���� �ɍѼR�2�Ve}�ԥs��H:��B���B�;�_�W�Dk7��D���o2�j|	���s�n���-\̉�"��^5�@y��*����-PJ���d��(�H�N-� 4���#�q�W�H���H=x��|�g<���{� эl=� �!(+LE�V�f/�5{�����A�2q�S&���l%�Q�#�H�PSM���	ͺ:���b�o7N��
�#��~e�Q�ۮ����?dr(p&
��`'�~��v�|������R��S+�-G��ǀ!\��BX��ϥꓹp����c0��lXlxV64EB    38f5     c808��8�Ĝ*ӑ>B��0
}�GO�P�8�uj���	�[(9ut����K���ad?��ڟ�j�.ʔ�-�۪p��ߑ2��<P�2HʆP�bRT�ҏ���������>�zoӬ���=�\�5ן~�0��i�Dɰ!���#��k��a�Eࠢ�U�tjF��>�6�caa��V	�ނ ��*,��/`�Ԓ����[DѺ�Xj@X�Tro�޹�%,�>��~�u�=������@�W��Jbe���ʬ��=.��~u���5�/��FF:����8�J�:'n��O�L�}oj��?w��͖��3wpXՄ��W/�bU�'�eqg0,˕�'^u��o8E����.`�#�~�2��r'|]���@�.�M�Xn���%��Y�6�yP�Ր�q4N��/�t�����C��'Lm�� 	�����Zd�+���[�4��$�yp��4���:&U����P-�Gl/MX�&�g+�<�Ҝ#b�Zݿİr`�Ǝ+p��������嵿k�s!���P7>\�~]�y�K����bảv,Y��V^���e�#���?�ӌܾ]i6n�xDj�D�9g��&n�g�>G��a6OR�iK������+�ʩ,9�1$ClAp:�l���-�M ��yD��ԡ\ei��|�;*�uӎu7�����2?���������w��� 铟�@� �͖�r�Q������-������E�!��&�;�G�	(����_��'i�V�\ڼ'�,��K���i���bJ���������;�9sd	��{�+#ubdN����U�(Y()����Q�z�ھR�q�����J�S�����a{`�i�gn���n��P_� ;����X��b�i$����-�v�E�N4t"K���|o���!ar#Y�kA������1�+
��F��u�e��䤭4�!��C�2��bb�,B6�]����a���%~S�ϑ�yh�~��Н�Hɩy �pڎ��ժ�.D���Lr�_s��2�h�Rl�DK�G���ԢUKrm �-�''����99kc� d]��I,�]���E6,0����|x̖U߿�ܿ���能S咱Q���A	��MF�SO_��M��}'��S��"-���$���L吜��c��01��A �5��~}�F��13�a�X'ʛ9��^] 	�K4E��B����KU��Ju�ܢ�]I��m���Ih��L������&	~B<;׮ ����'{ 
�A�"�����"B����~�J���jV[��ڨ��黎��0G���b H.�u\�[q\�ʽ����}OK�'I[ϱ* ��.���6���j�RM�r�SIc-7k]ևl[�r�t�.�Y��Q�In�Ǚ���N�E/�D�Q�G׋)����t�Ғ���/��
G���i4(�/�W����vJ���(��"lBJ3i������?z�E�����-����;=�v�(�/|+P�M���D����L�&̥x��@�Ц� �*4��b�^�@$^@�XqĻ�����,�$��Ȯ��3�5.���'���DDV�����:� �栶6/��}���0v(��03m�����hf�M�^�o�Z��r:�X��Īz	�CT(x�w�anik_	h�XFd�H����I��}Ѹ�ÒRG!���������ĥy9$�*���_kb�&�%��v"%�Da�y#
LR��K�\���.��!�WFi��?u�����KB#�>�L]�eߏ �b:	~�ȑ�����ı°um$y�f��:7�ͱ�H���������Ҟ�����km�v� T�L��1��w�� .֕7���ulZ^�Չѯy ��"�#�pֻx��RD�v���񎷧:����<Bp��7�f�@Wv1�Ú��o�$�5B�mhP�R�)�G aȸC��L�S�'����N�4+�?e`���&���,O�K9hA��C:���L3A�je�;}
�߿�ęZ�pf��.o��oݵ�� �m��Y�I�2�����	�Yr����-�l������'v>����PH�����E�~���Yu��\�*�|!VAuv�Jp����h�B$C����1��e��يekK�\}��Z�&�����t����y`;,5�ǢK;���\�lT�F������OΪH{��S��ԣ�ǰ]��./�튠E6�)����t�d��(b�ݍ��(V��������jeΣ�=��0S0@�b⨣��%�d9���O�1#�ODr���#@p68�=<S��X������?(����<�1��b!�e[?G٧�-o�F4Se�ڲAX��%�ɷ�I��� ��|ns�
&��;��{J`�Z� �Q��ṿ��h�*0'o���ަS�(=�[t^�3�p�ofO�����u�����T�DW�e���=�ط�g��=M��������ʃu��c�pɖݱ
L�����`V��#?��6�k�m��	�.�C�c,��%������2m�㗧�mMۨ��������`�ux=1@F>*Me�oч�~#��
#�хN���q빬��?({1��(�6X� /��	R�hX�p@�Il�������20�r.=e�,�-["~G�|*���qB]�	�d��Ҋ��j��a��� �~,"ꈺ�j럒�G`3b�Fm?� �;m�L�0�^��[��3��ʍ6��;n���d�>y���/:�k5���U�1�MR�f�3,��t�`�ě��H�卟���⬱�5^�r���Js�
�lB�.��x�)��A��>o<x�5���cDp��/b����g�I��R{>p۾Z��gXJ��[�$��vPY����'����Sڣ��^zo�����΄Et��'�=q��dLlK���\ �j��#ʅ5|���o�\#���7dBr%���-`��?9{�G�Bf��,��e�+� �ԴŚ}�t�	9���}�C��|9�A���Ѐ���m��=�!J,�����s���#gTi�r� h��j����	3��.:�ڑ�.W?W%�vR�Ud'$k�2x,x����C�j�/��e��?1Y@ؔ��a��󏭞��G-xGTd�ߢ�C��/���ǂ׻8@ԎTh�b�