XlxV64EB    b734    1be0�J��:����C�$lQ�` �r�����G�M߫���U�7SU68+% ����2�-��&�?#X�Y�ď��ƒb���K�SZ��k�|�Q�#,�I쪑��F��q%��������ĕ���`?��vb|]!k��|:�
3�rb(�h�=q� �xF�4(�+H�uҫ���"XЊg���P�I<��X�:�7�mB\�8o�}��� �@��� o�G{�7NZ���!����"D����Q���b�����P�/�q�04av��y��Um}�����Ъ�?�@�YPd�r�������Y�L�
�ל���������Q [��W�Eľ�1��l��
��Z�ƻ[��[+D_��N��m�`�����Ƣ�Gm����բ-r�����5A=on���4��Q�o�.H�|�����e�Oyw��,������@�I3��P����y������LY"�s!��]�X�;'��\"۽pd�����g�zp&��k����θs��Y���@�;��� 9��wT�.��	��Z[�1Eޥ�UL ��O�69,n�<~b���3�th����^��=킥�U��H�z{�3@�돺����_R����#��R��\�>�j���J�����h��3�^��?}�y\`8�<��I�I���Y��u����Y]	�y�!��z�Ӹ�_=-�V!����hn.��"�G��_
>,P\H��;�xaݰ�춲��7l;X�Mb�1�~3"���4Ю�$��a�0H �Fasd�j�Ί�P�t����c���ӄ>���9q{�o���, '}U��}ȸ*��e��b>d�y�1V�����]���TzV�x��MB���5ҹ�T����=#�ݪ{d���MQV$ӄ�X+��"bN?Th>2T�.'D��}���`��j�n��ּ�P*��Ga�k����S-�H�d,��"��ߒ�,���6��+j��be���E�ߋZ �]��ɱZ�!�������E٬�SإE�V\�ͽr��L���E�n�8��1��M�LQ�&A9�PM�q�k��d��ͷ	��9꒲�PD�z:)BQ	#uZ����r!����j�������#��.>��w�q �y���� ����Lz6Y���,F�V�� i��+�1�[5��`��`00�6	�l�m��Z���^�E���)��#,UIٔ��x�^�*��n\r���=�N�G	 ��� G��y��
�ȠSM(�O��JLx#�}��~��}�Z~���wt`�ϥ+��@~�a�RUVә�X�N؍X����*��rV��o������o=4[�@μ�gK$A�Mwk�\���c���W��N��A�*������j�H�5���w�@F�e��C��N��m�;����jpır���-�j!9����+!JwG}���d�����ݒ1E�O��`b�O���x�8������mq�p70~���T~���C�:�$/���M\��u�c�����y?h��R�2�9F/��W5�\��/\|%�8{!��F�f�*�;���#,��%t��g�uG��E���]GU��0����|L�O����u�Fc�j�-4���#�N&�EB�t���y�uu�F�Q1���2��T��M�؎*ZqK�V�������tR�u�T6]7�(|���<���P�)��&�����0䆣��A4���,<�����v��ŕ�<��s�l�*�Ԉ4G��W�I����T�30�O����,����R����6{��7�����{`;��q�-�-�4S(��R�	Ǟ��0�Ŕ���IE�&�c+LS��xѹ�ߊ��JG��)B��8:I)�ZE� �NEK����$媾;�/q�����[l��s0�~l_�ՙw�.S��۴��yj�r������Z7�[A4�����?�%�hgo�C���!�����oFȫI�1����2���lot��y�i"�MY�R>�,1�~3�'���%a����gKG���rTl�����|��:���d�bl���km�f�W�-�Z�."�1��OuO3؁����DX���,�puP��^�2��>���1ā<��/QQ�����˝���/�?��O�њ�Y���z��(�q(�L��K,�Q�P� �Н �s��zn��A��і��nƂZ0��-�y�]������Y`�=V���f<����9F{�/�YHeA#��T���!/�񑵓1�#�Or�{|Z�G؀71���$@VGz?@���f2P��j}#��w:��+�HQ o� �8Rl�J9?x�z=�2���ܩ?��Q�V�l��p����3��>��*�2Ɵ	��sA*6XX ��T�#��J��î�,�2GZ�V� ����S&̃�_��R?�?��=�6���C�S���䓃rԜr�Or���q�q��*��{:n:���vY�gm�Y�.t��|�)�dƥw�u��cK[���O�?:}�71ڳ�CX�#A����z�1'�H�v�lg�֦!�p|ݨ��/��,����a�0���}c�Yx9F/�Y�B 8�1rn����T��):tJ���y�D�A��)�򐦫�A����)����}�o����}�7�D�$����%�a�A�
��]fBϹh��Ƌ�sB�>���ἱ��X�^[G�@+�l�B#;,G�y&8,<4�13������%���%"��(b�j22�\�AE��!���L5+Cu���HX�������$�O`���S�'�%'�8���IA�F��ԩ;��|��VBR<U��5@�H9� ���������Ȑ�%�<I�/c������=��uE���=̍��*�&E�֗�ݱ�O��r��Q>�;ǳ1q�M��^���w��2O`§�ƿ�a��|��Tuc��U�Bi^��8Ĉ�U���������PD�6d m���-٠joQF���$F�����]�k?�hɼ��TKXՇ!��GN������b�ڶ��|����%	�>�Ɣd���c�$��Z)������z��4sX�s�D.���ߓ��)W�m�T��)��L �8_��� V@����\ra	��,Ύ��e��k��=o
s����c�01|pw�f�#h�b�?=�p��PW��_����R[p\�꣍���à�e�l]�\)�1Ӕs��}��sǷ;��ڑ�KV��:/�v�7^5@�%����Y=腎�M�}������sh�6C��ǅQ���_`x ���e�h�l��i��LhG ���֛�϶!{�`���]17Q/�6��a��V����$�K �^REts�"F3�����bi+c�P=�@P�:���t�랊�Ygy���m��9G�%A
��sO��3������p�櫹��}w��]�[�{ ��k�)�su@j;ǆ�����~#ڣY��:ĥ��p�kCI�
P�MX��+���U���,�`�dјʍ����Ǚs�ٿG�l��bL��T�J$/������8_1\;�V׉��O�N�@nV{����?��y6�el�z�W���A:EK�c[@�ܱ�K��T��Twd�����R�]Η4�ɉ�A�=�r^��q�(?/﬩��<37��H�H�y�y
lj@I
M�/R�MiT�)6���3��ںu+sz��Gbܪvh�P��vg?��W��8�蠃_B/x����!!Y)0>R��V&�))����߻�GS�-Z߶��~��:�]F�<�63~z�݃�k���}�Y�X�wQL��bg����-�^�>�c�I���(�!
��a,ˏ#��麡ˤ4���Ԛ�ƃ��7G�-B������Th4�j�p��C�����c�gȢH�m� ����:�����k��'KSNr6@�՝^Ao�͔Pv0Y��l-��U�e�[U�e�jG��U��� X17j,Qpv��[lH����au��G[�1&�DL�-S�3Nso�e��tk�5=I�j;��F��b]�[Cfm�pk$1�C	���[���=2u8<e����-<�p!̠Ði�K�V,dbሂ���4�ǚ�K0��~�.�L�@K��!u�(}B�S"9�R$R���6��v�M��&VU֋So�û��x� ���s0U��~����+�_RĶ,�W�i뢛�Π6�x-��>����zo�h-UK"�6TQ^��=(8~Y9E�: 0R�41&ԫys~��ʄ�B��9�]��@.�-5�b�<�B��#^Z�W������\��J0A㿥ԭ���s���8|��'q�1���)�����h�H����,4A/�˝긽aw���d@v����[x����`�h7}^d�,5Oq������Q��F,$ȑť���ot;�K%T�X�b:bС;[�*e����Ʒ����	�;�M�����8
[��|��D��� �ۃ�@�;�͹q���L�[C��Dm?D�;�r���r�|ܺ^��@�!�3�7B;�[�7�>�U���c'�<ƒ&1z�x.��d�śv��j��|ɠ��?ݲ��ȯ�ϳ�h���^��&M� @��[��������S� ޮ��-�/�m���� 4��N�W����:cXǇ�ISV]�&�	*%`����Gu��]J�+�B:8%t;|���nY)���@@�/,M8���� i��o��&U���Z^E���oӫmaǄm?U���Ժ�-\�Dp[��g�g ��)U>ҍI!���$���N�T��h6�܂�f�+�}�Kx��}�1��fJ�/�鐜��j�Q��1��Q��I���͓)�xُ������oԺ�9xG|ɹϹ��ȥʙ�.��ʉ?�zyO��Q��+� +���s;*;��u��Ĳ�L<��WdqjU6��X;
�M����p�(e��q�![���E����r�~��&�9ݬd?�5�����
4(���UA-шV�M`��������Ǎ����%&	U��E�Qބ]��[����l��~fK��͹Q䝇X`hG�)d�^��3x�W�)��P0��R�� �m���$�v�E���G��8's_�,?֫�`UPM7Q��zܥ_��hGdJ����Ͱ����UD/�ݿ�-:�����^���-��/*�=e"�#ɮ�e��3��ڦX`��a�K�]Z���c�	��x�E	OA}�Ql �/ۍl@��N��Fs����5���\���9�x#[��l�dTu@�++|6{��N sGܫd�E���z�n���^��	�aM��<�S7�*&�� H��Qd��&�����Ҫ�̴c"ӊ�����Ѓx�jO�%��M��Ow�?Ʒ>��rP΃eK��k�/X�-r*ɒ���%�[Q!��d�Z�3���G�=�2��a�L�v�?��"��7㸁��B
�����4$�Z��ty�R��$X锚���a=ٟ�y�C��s��}�`��OS�p�����WR����ȤIҎ̸��TP�~�#��sr��0v�:�T7�����Z��I�Q����x���6��S�k��~��{�`���'��Q#���y������#�;�@��io6������;��K��ʑL�*��$i��{w��ۚ��dQyV,ܢlN���+ݶ�_����TfV����n`\!�&5�J��A�=ĦA凉����|��RGR�xf�8��,>�\���l鯽yyQ�P�Y��,QSQ"�߆
��{��׃�iH�A�b�m�n2,�-���GZC�K~�t��E���c�=�G��\|쐩ݨ�y��pg�M�^���v�!�`�l}q��^nq�4�_Z\�Kc��?E��(F��f8֛�ߝ/�a�Ɯcfx��לdDU7���)��t8�w�0��j�wD��Y	�J�.�;�uN�%!�˜���uǘ�Ÿ;��e�u��4t�[[�;H�	zV�0��H���Ĥ��r��4e=dn7Q�l����ݨ�����ti�=�/�&4��tU��bG��Ǧ��bŝN߇vp�-�"�Tw���V#5�� ��.'B4�[Љ@�,ȼ��fJH\���F_�U6_���+�A`�Ҩ��W����BnS�N]q<����6��>'S3"��^�����@J	D�Ö��C�	_�k��ʬӘ���E�)曼f4�}.���J&�ّI�@�_�!Ι�:Z�����Q��e%��~��1(�M��2eX5h����/u��$�x�S�;��->��H�����R���u���4�-�ט3Ԓ�3��ܘ�* �<#1u������~���ACр��
m=�S"q����4a2$r�C��4ݮF�Y��`��[��������'	-�>ei��ː`9e�J��tB�X�����,��}�g����,�2;p�bbm�/��D��T���7��㼘$Y�e�~M1�ǘ�܂�%��U$����`o=8�n��ob2�s���H�2}Z���TK�,��{"�\֗LQa�8å�ܣ�A��2֕+�����J��Žw,��-W��P�4N�V�@FJH;��!j^�C����HH�4�:�"~��]4�xC�ř����0v¾~"5��Z�b�B�zZ�>o��)_n� ߖ��u��}��mr�L#�T�T발y���=W�W&�ͪ��	_L�=�^h{g�r�f�S�C�!I��M��G�{��ʞ[i�ծ�p�Q=����03�_}8HP��Bȫ ��W?pn��3.M���D�L�1]���i+�J�Gm�r�{���#����)l8��rH1�
)��G΀�8��������~;7��\Ѷ�ت�U�'�>nH�^���#Pw�c�ɉ�M܍����au�xy��EEh};
�s��1*���:�gM�Ԁ�{���>!��G�fP�����S�R�d
�Zi�J��(25 �л&���D�~�(rfF�ηh�u����Tk�y!�w������:&��� ���Cp�bH�*}LH8��}��l�C�Mk?��bN�ӄ�ZH�`�S��BD�dЬn����7�jT�#3�ʓ���*�'&�xd<r/��W?�#�C�,W��*����3�X}�|s�xzF���N'