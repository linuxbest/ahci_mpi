XlxV64EB    1b7e     9c05��R�=H���@��K� C ɏ+YCi5�4&W���%N>SM�#�0�$��M�p@�!0(�˸/��0b��Vs �"T���S� ~�AG�{�̟vcèB]%���~�o�b$��<O�t@�_��Q��U�?W&��q�
���h"���I��S�!7�Ԝ�ڣ�9�I�@�LY�ht�է�|�+�|q,���5�G�OR���e������I��V����T���(�����=C(�յZ�q=e���Ⱦ��V�k�,�2H�BePʔ����Hs�
��4�T2�*�"�V��'����p���해#6򣚊���i��eO^t�`��B=�8���=�L���h�l�*r���`P�	����]�* � ������bH�!�4^Y6ԼE+ 瓩蔈Z����tQf�&���̹��,��y��:��7S����nW�ˇ�ٯ��󋚽����К���j�`Z�$$�m�Z6��Bu�;Q��c�.�<�xe�2y���M�T�E�������^�vc!�薛�9�,�bz��8�F��S�ѥ+��X��!�� �0O�}�Њ�@[�.(�,�]4J�D�&�:�Y��^��"��R&Qn��W���cx�o���8K�����ݷ�:\�y1.g;��^�Y#[��b�rW���?t }bD�f�B��@ܖ���5B�����/���/�Q�K�Vfv�d�y��U�jTu	
kG� 0�i7Ѡ�
v��)a�Y\�\9u��~��>����$,Cg�@Ғ�	t�BX������~U���Г� C��q���g~3�Z���~⇐��}�I�/�������s*�A�eëbz	���M��ö,�'XԺ2qߪ�w�X"���Rd�>��׵�Xe���%i$#��O|mJ��R��s���V��q�� ��,�8�P��b2k�:w�?6�kW�:bKUA�V+��x�ķ�	
�<�$|AF>��ָ�7�"�Sc0,�����↿��� @�u�X3�[/,0���T�n��Z6B�<,l�(������@�G��6È��3�Z�s�<�E �`����Jr(�נZ�Z�(��D�Jx\��g���I��(��
1H؂�ٓ�~"f�K]��I&@#�s��єG�!���Cφ��W�@����|�.��Nv�jp������%��B��[�I�2�w(�_'g�CSp���!�e+8����p���W��Fc�c���#�Xb'_�e�G�Twbn�a�͘ң�ĝ)�i���#g�k�9��\GO��4�s
�Hl	v�Xm��KI�"\}hD��\~^���F����O��/���3��4�@+ֱ��^��+�|�}�����:/h[W3M���zģIѡcn�>*��j��P�z�"��A*��D	�J6��]�x�t�^��[I1�c>�QK�Ʒp�7�AhW�n�-��b2�`���#ϼPw�5#w 8����K��'<�v�h��^���n3?�!���Kֆ;��{9-�F����SMY ����g�C�C^3�3#�j�!�����H��
� I(��	Ϡ���(oS�3��dY�yנ�^t�`��ē�[�K=���3���'����R+'R
�.��K�H��6ݛ��SJ�]���W����Z\���b��p`J	�A�����b�����Rm�H��f.��"�{� nw>$V�'@���@X�ců��)FIacw��fM���,�=�ey�	'P��>�e��8Ⱥ������BXIX�����c/�n�R���p�u��AՏܽb�5
��MU��*�-U7/�h�Ύc�!K5�ҕ�����?L(�]qC����� �蔼E:�O]<���u��ϫv�U�YE�9=@<Jq-�4���1���RXh[�ɟ\L��d�h7!H����-��	�U0�6d3�x��&.��\�mnΔ0�Ό�57Yi���tӭ����\��F�-,�ZՕ��~d����/�ʂ�n�!ϒ���YBC?J����|��NQ<�=��,"��n���C�x��7�+��z�ap��� ����^/�����3z��ҹ��eZ�-�7��l�Q,���M9P�]aB^����<�#Y���r%����Sh�	DݑT���O��>��*��w/�aC��x�.��G*�X�q23ըPt� -�&��K���%M'u{VnkL�p5�7�o���o�=�Q��67���:>�<����9�0+GU3�ze���T9~tG�8��g�hB��e��u�Ȏ��_r�C>/*��ʟ��
�P|�0�>Xj`_~%����|�K6�&�5
��v��p��������zA30Ļ�KQ����`�.�șqovR��Z�b�MR���a�@�:$~��f���(�OoȳZ�-�.���ưDR�F�?__p����O:�|� v۴8��L��Q���,%��|5� ��-�<~FQ�Ϋz�U��2�^��V�2⛢_��Z���