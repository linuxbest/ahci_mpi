XlxV64EB    48c1    1290���P��բa�
������߭��6 ���׀K	i[
���SN��B�U9ǌ�]Z�=bYү�w�����~���4d��Կgx�D�Mh�jEΚ|<��\A.X�C"��@Cc�q���mY{��+���aP�g�*�d�i�t��5��.g��y'����i��Y��},e��-*G�-��ɸe(�Y�7��O��By�p���&�qdSH�����
�\��IB���||���K�Pʛ�'%T���B0�e�.���~@oG�Ѽ���ۚ�O[��o�#�n�sM͖ER)8��W�EQ���#H*1��u] �W��ƃ<앉#Y��!s�����;C���u�5!�p�Y����2��
�@O�9�O���JM7�%��� :?F�㊆�V�-�>�6�3r;cϹ�&�nZ|"��9�u�'=%L�Zډ�p�I(E�R[w0[аR)�����aLi_�{��1^����s�S+�f�5.k������~��%��Sn��3ߊt�Vu�i�}��=������=m������[�W9����7����ei�Wbi�g;�
�����;1�5:ڣ>IpⰙC&���O 4b���0��C?����H��duc ��3�Gh3 mu(ɕ�t��8���-Ą�$ڢo����}�$��L�~��������Е��������~�Q/��~N)��Y��\����Z���R��S�֕�S=ײx����jK���J7M6�.�yz�a�t��g��̈́��H��\��&���M+�莳�����!'e-6�����^��$'T�l������0�0y��2\$q����?��ЇM����.�����o��4ތ��1����Z������kЀ�T�dl	�@���%���-��`�M�C6��-sy<�$���b�����vIվqk��l�t?�i�5yb�z��;0M�/q�Y��a5���"�l�t�?���<�S����ŧa���-)e`�p�D5�����~2v���游xC�-� �
!��ˠ����H(� ���r�e�-�p��o�GG.K�p+6��\(pM�7����f�$OέK�d��L�Fƈ�rwGó8��RcW�v�9;dV|�[��=�o���8� �{�J�.G���[�����tK�M��,��#b6(�@J����f� �~���рBEm�2@9ʊZx�8k�_$�"�?ӹ�{��q�l<r��/]��c��ǡ�̎�����������}���h�XB]�"��,�����(Q���E�=�z=NtM�T8�	9�&�	�O��!33��(Q^\�uq�%���e�Ó�#�0,�D��y���Eߏ�0/��a���Js5���f�%����^e��^���m�����.���灈�Ĥ���^J�)�^����7y7��7��*\������[�B����zJԡF�q��A��"����=��N��{|�(���x�~6�.���E��/=O6��Y:�����p~Yi�R"@�tg��,����"?=7\�j6���2��7��� %�*��b�^K�z5;wP����
�h�U�L��4�}�b@�?EY$��?F�/�C'� �Q��<�}F� �Tx�%5`�5�&��v}�c˪ц�^�v�g�����ǠB!�_�\���ʬ�1º��(������!�����F��^͗x����S�Dm�`E<�u�zG��׿�Zw޷�
'�A��G��n�׌���g���B����r	����8�O2g%�O�p.3�s%����Sr�K_�WB��]`���H��u��0f����}.��q��p�b�^(���F��+s�>�u��TRr)���yRv�z�crNz��7m9���6��ii��	&Y����O�|���G��P�����%���� ��b^�X="v[8�[�R7�y��ˀ4�3I�Ք�g��6&KiL�M���b1CO�[��s��zya��-�ؕ���x���aM~�4�A@���۱�騱��f����1�2}��cC��MJ=DNh���E
����k�`Q#�k��z�ıӁ� ���Φ��O¥�����
��)�!5r���y���-��3n��k����W>JJ%+h�ƿ��zm�橿��ֺ��:MXjNQ��?p��~~�[��W}Eä��}�y��k~���^�3!Q����u��M��F�� �5��-�ZW������s2�L��i��.�,��K�a*��D��l9��r����t�����SWRo�I*0z8�!׆=d�̶	��M;��bLn��̷�by#������%3�Ź�ID{%�X�Z����h�R��xχ�C�K�I��� �TǄ��@=��ማE �TWrTR���9���iyN9K+�1�H�{��C��ŊlN#@ֹ1<��"�\�o�>S�<[�BQ�s����G�:n�4�Z��ߺ�d��I7�Ω�7�(^���hjO@r���C����xDD���i󨑃����ǈ�I=���'vqr܇Z+�Ԭ�ݍ��R=HGt�[�'~�"��l�i����8@(0 �[i,��R�R���GUݎ��,J�
- �S�Ht�\Q[ё��Y sSj��5{z��?�
�y�2@K�藝y�=C+l�����7W���Z�)�֌�� vͻ|�r�y�i�gj�}'��N�i�$�>���s�<J�bP	�0�̆�H3�b+S�����y���-���3��3m>#u�E
��^���{��g������e��K_R���_mb��t�>��g��A ���z�%�T�c _Ak(�eiq�I�󉹧��݄�%KyJ����ml)y��&!=ZK�?�{��m�����uW���N��j���b�ߩ�G���i�&���d�x�!�e�42���|��6�d����ݺڷ��-Y�!�m���Z\�wV;�(���/&H[��;g��Zab<@`�`w�jLM����'�N��W��g�(�F��&���H'?�t�1��S&����p;NSD��غ�M���7_q�@p���FX �Yk�N'���9/�S&��P~�'��]�JAW`����CiFݕ�l'�3��;�K)VPF%�t�f���l�T�jy^Ή����Q��-��.$ݹ{0o?�7c�+d���:Ű=6�~�����e�N���I�=��E�k�%ܰ��
�vA�J\&��%�V�ئ2�$^�b8�K5�je����QW�3��R����,�y(n]'R�m��O7$��:�F��@d�n��1|S�F߾�a�!lY+�|�"HAw���@9\Pe��HĦsO��(��\:���!4P�����~��w�́f`Sz���������\����{L��є2D��Rv"�o�X���0j�P�	Nrk�'&%��L芺�;)���!��N��9eX�w��7��"�"���Jʡ��-��3��ш�)A�RpW�@�?�fyFs;��XQ������`{�
�(ވ�����]�+6� nm��l/��䭞�7j�:ԓ4׉n�B_A^	%�͘Fz�*���vwY:];DfK�0|��]dv r����Z���w4x�J���_���ZV���$z9�����ʩsZ��oF�"�\�S)�(l�d"�/(h�'���8ǉ��M� ��s����Ku���Y�	��p����A�Q����c:���f��ivFphbD�qS�z2�aP���6���.�]�xx�T�X�I��F5Q���UC?�q"�A�� !y����^��e2K��}�Ҟ��Z�pI��s�!� ��6���g[���ǒ�Z\��23@E�gUo�x�.�:Z�!�����d�˜a���AɺB�AA�_��=��f�j5Ç`�pl��]��!Io3巁
)�C/��g���#�8s.�q�����D�����o�l�mq�uD���<וQL� �slz�o�|�y�Ql�����z�5=�E]k�Te[5����?��e=��w��\�nh1aĎ�O������ p6*�~�w�2������)X�w���X�ؒ,�iA���������O���N�;*�4{�>8q-��A���βd�A���/5A�S6�j�5%4�R���Eq����C �~�lz˨ Ml�������_�=2�;,h����L���X�K�#/l��R�ڿ�������$>H
��/�*K`4��`H���g�!������ɿr������Ա����T�!u���Z�T�@c=�}Hӆ�f����k��L+V����Z'2�ņ/K��e�Ѕ%䖿���K�h�Tg^Z�j�X+Vs��n Z�{�,�w+X���.#��/.�Ɏ���@�����]$mh����&8��@'�r?ٽ�cZ�iy�jɆp+8��.߹r)-�ړ�ĕ��A�k��wC���2Fq.�8��%�,��_�,�oZ�K[ڔ�.�3�tA��&А��<M�.����J�q&��H6�L�U�B��E�ڛ�07KX
��)����_������G�9�J�b��c�xt��?`z�ж����ʹ��Դ��~�pjּ1��o=�Ly"����Qq �߮�]ȷ�e���Nb�{��d7�q�[�.�z�F䜟�Rx�@�R�����-�G]�J��L
]ґ�C��� ��u��C�d�_�c[��;�&ّȃ\>�