XlxV64EB    1f8c     ab0��eQ(1�4]7�r��_@!c��\|?�����`���&��Ai���1�[D��R�C{q�=�Sq�1Q�O�tT��¼� �nz�B�\�X���'k0�0��_kx'l�4n=�P��ŷRǄ���oa��Vd�y��Z�S�O5L;�s_}�Q�����UR��AGw)"HĴ�߿>�I F�E���^ٹrd�r�1j��Z���0��J/|�2'��Gи;�ѻ�m��p\k7�v� �0��ksVW/P��;�3ˑ~[7��@^�b� �1�v!��9�b�������Xl��]�gي�:僉�����>{ֵ���/#ǐCY�Z�ok�>zl_�'����G�@���%�^bդI7\zB�^��͢������M�E��z:�W X�v�,�"�G�s'h'mE�r��Ha'�d>��Y_�~�;O_���f�ͳl���=�	$��+�
�  =nB�ez��5�+L�Th�Eqj�cC$�u�zk�B9��W:s�א>��� :�ܰ$������3���I"J�x�gSoe��I�v�ȍ���g�
6� ������6籞 2gKsV>�t�t� �ݯs ���q���G�x�p@�8Ǜ穵���Ȃ��� j���1.Pq�@���(�.�e���jP}0Z�|�>7��)'�}2䣁w/��f�~m��]�P�� A}��O�p)\-�,��nt���&U��^���G�S*S#b���x�֗�afA��f��ʄs�8�i��:�H8y��?��Af733)n`&�oaջX ���NW�#a����\Gt E'�2�SVEJQ��3�ʼ����T�FM�t�!V��������ʘ�����]�K�jg���U��
�m����h):�Yz����?5~$	w��(Z�4�mAf.S>��$����N�1Q�'�̓k)�T��G�����ޙP%t�+�V[Ѱ(�˩9C�_��sr��`�Q�[�
��6r�-{������|9$�W\L�Y�y��dO�y[4�r�l�,�����9�:<΍?Аw�9���A因�X[�~��TP���`g8?�i�]��6�/��lh��%��*�,��:N��� �x9>'i�gr9����8͆r�|>5���)�;��Ĕ����x�% Ɣ��Kwέ��RZlM�F!�w1�m�ͨ����3�u@�sv�h�D0ϡ�Hf�!��U"�\���W	�U����}uGz9ǞWx@^���fv��t�r ���a�f�T�t�N��^�x��i��&�.m��H㓈
�'��.�S���1
ɫ�b�4j}����VR�͓<Ó�X���hy����ؓf�幣|rSՎ�x�tI�x���e���(���D����O��l6O�u�1�<ƀ@�ͪB�q�;_[&�My��"��袐����#R��\R�Cf� st��`�<��6.�d:��� �B�;�3�S��X[�O!�V|�H��tFn�n��?���1����=��c�A|+�6c�Ȁ�`��M�l�H���R]�p`���y��2N�6� �ݵ��Nd�@TO�t㿄�(3��5]S���H�\IY�p
�4��LntZ�|Y���B�zL�,?�H���xH;������ת?Z'~'��^z�)���+��}�.Q�ϳ�akG���Q��\b�,0��GK:��%�:O{��ʁKɒ����R8-���d7Z���lD�Ȅ/oԏ���YK��.��]�+=f�~��1o�
HѬa�W �ߚ�t��|����z�>�Zc����p\��w���t��:�K�׼���]���R��;`ad;�Z�5�
Y�ޤ��2(u���ג�>���Cm]t��n�v�$�S#��,@~��
����Ef)�u�\A�z�'S;�p�3	9���v�N�a��E��"UË_���;�?����Uֱ�\8P��#�v�2���aN�\��I� Rt�ܟ�:!㠯#�{��~i���Rl4	}�O
׋��=ZNF?7�L�ZX�c��C�ɚU���"�o��s��s=�+�G�$�fy�&
&�6,'��=Y&�K�=����s�Q��ɱ@�E��M�y:�:�yBX��2�ck�W��)%=�Ǧ	�!����-ׯ�A��ɴۜ, �[Ll^�]{xH�ɯ&됗��^��ԉ]�YK4&ЊMvھe���;�1j�3"'�U�c�~��q��Auԓ�������E�k0s����/�[zsN������	��tz�_��&���	�u�M�5���yiO��	��e���$�!��}�A=d��3��܏�F��]�C^�������u�,Y���Ed+q�d�z_����Se^��5$���բ�4�����ͫ�7ǴlU8-��$0�n��'Ѧ	����lJT_�����B�!7~�A;�,�o�1,Õb�uս�{ճ��� o7�*ni��Q��~��1ҋl/�����yP����#�
c:4��-�3�]{�ߤ#�P�꦳ :��4�.[�A{��YC]q��Ʀ�3�q��#4�k��oP��c��0���nz-���\EjOZ�� ���g"n��`c����*U�i; *-��;�so�7}����(�N��}��S0!�w3�ݺX���s(���H:�Yޣy{s�&�=�_2�.h ���"�ͻ�ɳs�ܖjs�җ��Nl��@$����8��ާ.�k��(