XlxV64EB    fa00    1ec0�:���@a�0����b��v�my�ڵ����'���e�J"abZ�1��gSdN0�bre�f� �����b̷���R�H/	^c�U��7�p7$��Z�������DR��M,�Ȥ�f��	ڑ�<7$�࠿x���K��]u�:c��^J>	��"m�X�5	���w�U��𿌳p�"Kk��Ű_6�l�l��\��bo�zs�?׀5��
ǶgJn�;o�)�����m�!>��rx�fjP�ȱ�s@��r�S����*�rɮq�S�:,[�o�'�̫�<�.a4$�(��@qY�Ir���{_�K���G�t���.���3����t}��~��{�
)�����
�!�y#0�M�oC
�+�ڻ�jk�yp�p�ň�6J%��}uê�q;%r�i�[��g�)��v�l"�X�ި��EC����f�4�]�<}����-tr�!%�CI뎛9���SDVWw@�c�H�s D�i*�ZyM@��к���gI��lXx^M��}��d���	%0��t7��)�$t*���`mE��B��4l�d#"ֵ��%0u�/��U7!?��7��%�t�>�70�AW|C� �Z;�E�H��`��hY'y6�,A(oT�YgM9�Lc�|Z]ϟ
Gc_}ɍ$�Y8S3O��ߍW��YtFlf6�bU�_w��ݘNH�6��zI2��������fQ���PY�[{*�N�]�_A�m����3��)A8��:+2 l
���%jL�,�Q�9K��>T��0�����]^hH�[{�&���N�LM�`نX{u��)Cl2���h�zP�e�>�
�#�ߥ���Z�G��q��+�)`ao�G��k>������Q`�w���[.ui�X	�=��/��Q��/�����x�U%��,mH�����0����}�,�����.A��p�i%���1N$_[D��Z���<^f�0 l�I�⋏�J��M�Ƚ5����{?��}����sYyt���	�	�)�CI���(��$���8Q���N�^if۝�y�u����k|�>2U��;v�:��b/�tr܋��%�0_Mp$�S�,r�
��q�5�\M���H�#w�������@�"�~��P���5�<:��VcA�;yN��o�7���)�H+�����݇X׮'�y�Ч�؜Գ|���7��(�_i̝����h<a�Q9{̾A"V�v����P��Q��b��?�3�lSy���� ��g3B����ƅԬUǿ ��^��&V��	rW��::N�}g+/"ڳ�E������+�C�J~3~�I��(V/�nY��*�Ʌ��;��R;�.u(��~ v�dm�w��������d���'����Z�|�h��.V�j`��J���MC�<!��۸����t���(�o��aiԢ3{e�J�(M$%Џq��)�R���?�s���qo_���g� n(�`,�EBt�a`�������MC]^Q�I_`�qJ%��7$�y�*�e/R��,D�`�?9�����-��͎���������z%Xǲ��h\Ue�}x	��<�J�Z:�^����쩇��(�u�=�H���P�8}*�s���<B�N�༕0z��=O����J1�K3���h\H�F�sW�W6avBڝ��K������IS�H^���{��t�у]$��v��|ӾM5�X��ikz�,���1f��t(ޮ��K��5�O\ 6�{|��C��H^F�&�G�8&T�yɁ��6|~�eE�yv
�Ѕw�D�չ�N브ASF�v3��M��[b�ޡ����߾��_�~�B�|8_�K�����f�+�հ>B��Kۦ��@�\��hQ�5F�i|ψ��|,�k��<ARB;����r�ݛ�W�^��m��~JK*�c��p��+O��=�,�ԝD�: )CE����#,�F�xZ��R7��$��A�I�b5��[��9�El�٨�?�D͒�,�aT�tTg̹�v"��O%�"�6�IG�$d������1�������
A�_}/�=/�]���ՌdS#i�x���Q�;�M��׉���xHW<s��G,�7$�d��a�v���
`�_-���wˉ��rb�U_�m���TD��-��!��	�Ǖ��b�#�bn<S@��xu�6�L�6��hp���~���ї�� 
X(�� {$�`��� ��4���W��Z�cc��q�*�q=�N��$����2�W�hc�����hF���,�sSdkO����Tm�s�
�s6qt��!���Ro҈���<��E���0�eho�V<V܂������[��q<>W@\����^>VO=X�]�l
�4[���:�Z`�|/�י
�9ԭu�g���&������ �=�/{p�1lP��8�#��3*��
������)�k����+K+$��Ǎ=ݱ  �Z��i�%	���ÎQ#��T�&?q�>%p�.�N���}O��m�lk� pͩ��2�
�v��R�9$�Nt������������i�~��JP�꼈t$D��C���o�e���kq�4�X�I!���|:�rz���?U���&k�.˟�HK3"��Z���D���O��=&���ʣX�$:8�+z�~���<���L��zW���V/����땭}Y旑 �WsNAF��6�%L����։$ؘ�.5L�	�ێs��l����uw�e�4&?#��r1կ��E���,��7';���&M�`�(-lI�t�D�T<q���J ���/�����y0�C-�$V������ īud����O��͈��(�ke�D~ p������#]Tm����&3��<�\���6��ww�jԝ��f���=�F��>�׃	�G�;
>$����1��Y� �~O9S�0}��!�=pFZS�� }�y��\��-��6�i!�4ߋ@��T �iσ�zL�̳*!~���Q�~�T�� r6!4|	`��{�'][���4��\6'gn�W���Oء;�O�V�5����<�� Q:	����ӗ������#���5��=a����i�����`�\گ����>O~�@�dO�5�%+��*�@�CQѩH�O�:?�h��ɍY��i{��+i�ʐmx�֊��.G�Ga2�z�<�z(A��|>
������8�lM5��a�<'�lnk�(�І��8��zS|��3�C�־o����.E+�Nk�e�.���T%�{V�i�[�.K����>�6���Y�2lS�����I��1%v:W*��剈� 9�_ɄK	>s��#���n�<�`o �AhYwY�k8���p�GϜ�Ő�H�ͫL�n��y���;��M,ȯ�R]��dӛ���G��t ��io����ț,���`�n����H�{��u{��ܒ	S�yR��HP*B|�����O��6�֌;�`oqs��#�
�159m#�ӆ(aY� T�7=)Ym}�=�Y�ʆY��
���� �(�ťkYD��L\�l�f�:�%~���)Z �)P�w�13��;�G�!�a�
'	��ȅW��q��7�lC����K��J�;a��<��BuֹbAw5�\�Q����%�e=�F���K�d�Y!#�	-��,��Ϣ�ӌα_�>Z��2�6�����=���.�)��kFJ�j%�t&�jHb��Ƅ��9��cc]zY �Z�[}*c�}D����������}�C�48 ���jm6�p !��̖�LJfP�t�K 	��j�W5��U������(.�8�麫�&�����\�0Mq����]�
�ݿ�-� �RZ��Ș�k0�HD?�ʎ��D��/�-�� pf1.�rRtf|̡�;B��e� BE���+7I'M;;��NX��\��I���.�@��}��&�V",�,���M��>��Swi*��V�G���\��}�@ &.��6�Or"Uy�#jB+�I~yc2�t�ϝ����B�2o�tZ�޼%��m˹�hG< �dgbЦ�S��� ���v�G����*cQ<�]��o��>=�xP�>�-���q�����iB�L�i.��{K�;���hMf�<	r��������k�ʋ�n��� \ �o>4uC,P���KZZ�xU���'R䇕>�pB �|��,�y���pO�cL�%:�U���M��r �n796�F����������i����6���i����2�UO��.�?���{�"A����,I��Mnq������k�:��� N�2 {H�y�1�.n�4ñ�=3��$�n��;�����S=�R�1����J"���!����n/Gqig�lu��K�b�,Q�P�I��o�Sch�٥�����_�܁F�y��<���Zp�*F&�lX�$q�ڨQ�U��fU���ǘH����yыt�X`��>�]�c�׌��T�;��+�-�m­@���ІP�+��JZu֞�6h�J/�0�2�D���cjo>m��Lz�M�r�a�p�t��^��!���:�7TLr��S샼��5"�^��L�64d��OՏ2l*و��M���i���R��}��mb����5Q��P�����J5Vl�m���aw]VRg?�v�?�t��V���Xq 
;� �xF������Me���:B���,4�ǰJ+V���̶2�"Z�N{��M����UԊ��':9��Zf��<x)d�*��NW��q%��,�Z� ;	��S�Q�FM��m�5�m*�6���U�%�vY�����R"��2-�G��/9wc7�r����� �$tҌ9���^L�~6�Mdy\k�C宩Ob�.�!>?� �U����s�UOs�f55��R�_~D�Ų
��{L%�>G��,_��+��� ���)�A?}���������N3
���'�^�P��Q���#��}&Q}@
Ӫ8xb�]����C0ЇQ�{�뿒�h�ɒ�gV�	KV>����ٛ��~	�_�k���r	���c.$�Z
َ��k�0% +X�T�p��~��D�K�[�J���vmk��];ަ�ڨd��D|R�&܅�Y�X8�����Ro:�-K��dUZі�G��-����Ϗ����9S\n^{]�ۛwO[l�������$��+Cg����}.X$�8A��[����[η�t*�0ZOӘ��2q{з�ܿ�L}�m�k#F���AV"����-8*+�:�ZSZ��e��qX����&*A��-���og�u&+�c�io��S���ۇ����J��=U&Ǣ��@Rs���
g�(��V�Q~���+�)�N�|�5FF-��}�������s���8��I�M�߆Gϕ�\��!��Fb��'9k���3s,ǡLA� ���I�`�`㙸�g���(]��{C��oࡰ:���\R(�?���Ӵ�@)݁Q�B����-�-vYY'7����[�8����Ïp�H�Fzh�5��"/QtN�-'�K�Y�Jd�܋i,ݔz
�'�Yz_=�(��WmB��
P���i� Ѭ���$�R�+{F�@&�,��[X�vs:/5w
���;�X�����B�\Ǫ�:��]��y�߾�:i�Ր�㛾c2��1J������L���H�����.Zv�1�N0o�����+��V�ֺ��_�5Ņb���Z+�n�<|4�}<������,�ye��΋H(D[��8���Q�Y�d`�[��+c�ݳ%Pѿ��5�����fʸ� �9���^c���㯋��mM�T@��������#�Qg�=��`(	�_�r9�G�S��?21�	��&�?��$�j�N��?C�-\��.�C��	���=`�-�E)��%�	c��yj�iu���2\�U�]�K�q��6>�W�/ @����4��h���4z�R-��?�q	R�*�Lex
$�j�9�p_�r�:<o����@��9�Q�к�@t�t��]�J�,b_�AL&JU�1��F��|0}f]0=�����hL_i8�Ku��>>ZS=ӆ�i~����Ʋ_UGMM)�0R{�dO�����Hõ��'TY��D=X��T�#�����ǽ�j�t�Fc� �.��Z��i���B�Ϛ��f1���_�:�衩l��"|��ԸY����&��z���ω�Ȭ�[�g�Ay�0���e팪:hZ\��d��H�a�lK�9�	n%�����|r���w����m�fc,f�l��s����έ�!gdb�U=KZ����m��*R�_n;��[\�����
�\�E�f)�J��}NV�Iko�o���֝r����5�Y-2<aл�� %�=�UC��]pVf�A�\���/+�f���#��k�.�_�r@�v� ��'�ǟrO8SH���n_�X!��`ڕ��5/���u8pQL�X$}�
 k�� |�9�޾�ץ���sr:��?�b&��g{2К.J-]�	�7��M���q��_t�����Hz����PaoJ@u6��I�Y��������q���s_wa��5��c����:E�I֕ĭ��dn>�2/�����	av��Ǚ�� �K�;x�an�-t��>�?��Y{�������-p�����2��h�Q��֏En��-�c$5ĭ�dpC�!	i����X�`�6\�s@�e�,��lX}*�FQpdX�k� ^�E�_(߳���af���ߑ��2���=���|.+�n{���v��:�U��ObF;��V�E}����%ah����Α����@l�qU�B2�#FXR\<>�:8*0�<n*�V��{|������r��$��j����ȔxuB��V�1�{����9�5s-#�f��dj��c��D��W�͸z�T�+��;��z�]�c6�4����$���q0��|�3|���Q�}�ʹP��H'�g� �C�b�Ne����>�z��I��H��D���T%e���66�=|� ��5M.�1����������'I�T�F4��r؝�1�M�G�1U��5<ۮck��|#p�2�:M%���߅����@����w �*�Ұ�-��(��!o��T��$D����Gl��器���d�x����}u7,���f��2�D��-n ���Q J�_��x�Ͻ�~��� �=��V�
�y$�(v#�6 󷕌���!}���9������{q���G���Ѿs�:0Ж�,�k���������b���	��B��"F/��Vΰ��L(&61��g ����m2s��ݯ��"DB<�x�	~�9�Nõ��C��7'�u*���N%e�]����ЭU�e!_)�S�N��N��F�`v5���N�Eś���o�@M����L�pE�Q።3�S�g���[<��aVE�B�D��qew��T1$_���S�V,�Y��c̓�ʚ�I�DE>�$}f�u�O��{�)�̦-i-x���Jf�vB����VѲH�����G�׀^�榛�o���I��Ɋ4LcGN���Na¥���z&�{�a�M$h��g��{�
���&�Y*��zH�f�o�s�(-+̓=����߬��C*��WYu���`�H`a)2�3_��/|'�	���9������<6�gs<
#��Y׎K�����N<��-H�FI:�8�(**NS�?�e?hH�DЭ�|g�ltp�,�O<�#������i<$֚
�� �v�5t�4�K�:bdB��o�'���w�� w�V)��269�S�˗�ۭ���0��@�����
�A7V�0��OM�eY����b&�XlxV64EB    7be2     cf0�:��VT�+星����dtW"�h���j��0��Rp��,�д�0��8��o/ҲrÇ��쬨5��V�Z(X���,%��c2��q`uuH2���g�:2����5-�(>��@��C⡈f�&�S�G)	mM��b9P�W�0ބbW��%��н*3l5�(�=�M�Y�{���?^ S�tI���Dt���q�,A��̂����AZxy�S>9�v.K�M��q|�^�K_��$o=��<��3����y+�����B�e�ڹ_\;��l�iO���=|;;U�np���O~�=��>`�|O�@ma�Bh����":"+�D�R pʋ����e����;��N�A(�D�ۯ糥=���|crS���]G�P�K�e���&if�Ѱ��t�Ӽp�EG�Z`Ӏ[�}��tQc�$5b,?�UZ��z�J�+꺎Z�-�Ikh��_����u,K��Uv�|��ʒ
���W��0f�����B��@�r�x �J���=��	#'��[`�$|O'�_��{��?Uȧ.q��ܸ�l��!6����6�)m
+
���1�|KnD��&G�q!6q5��B�H��N�߷����ا�F;�o��	"O��8��׃�,!��T�5�R̬dl|��<�"ZGM�C�*�H�>e�p�sy.���}D�˝8P8����mm�*H���k�� &
�KA��d�E�Dc�J�X�Y&�A���%�O�	�E�䇜�M�5C�20�������24e��F&���&W��D5c��^Θ���֫Os�l�Ak��#&� Y_(��2,��ex�lCJ7u�8u(��y�`&�v��lN��S�c .W}�Q��N�C��֙{ga[�Q��`�߲�?o8�����饲��U[�A=�	A���˺���A��ſN���]��|�a:?��/�X�°Kl������.���%��詳9n�]��F/�o�[=U
��(&��=(@�^zr���Iu�}��ss^�o�<��\6A�������φ�L,��3�?"�,����Ttl/�� [e�	�'�v���8���e��$���2եy�o��1�k�NQ8�K����9�B��s��%jKv�g:9�z{L�.�7�:;�⪞�;�y$|��˪G��_I{���@�'���Q�3�S�Z���X}$���n�h�H1���,���p�\��ө��"	��a�x���WAή�m�e�x�uٌ,���maǥ�)dv�,c@	wZ���*�3��v�$�`l�w[��]���SkQ"~$><Q)�-������Ac�12R~���_�|�X�I�S�g�*�SGl�\��p�i���m�� �,
J�Є4��mI�ֹ��6�=��Fd��{ٹy����+l
��TP��Xft�zF}A[�|� ~�?�������7��ZF'�Y'�p��������n^���P&xy��*ǔ0��@Ɵ2�Z�~�D���z5��>�sd�U}�p�\���x0�;(������Q'q�}�TJ�zG�Ê�A���PCR�*T�c� ��%��^����u����>W{@H��$3r`7��X���!�-R�L��	H�d.��j]��P��q�x�/b����h�Vb6^<�x�І~�w�����?zk���F|r�g�`�vkՅي�=-$[�P�c{W,JV�RM���?E��پ�`�-,�}�=�0hq#*�t�wghs�C�f�OK�'�Ug�����F���-g��O��9#"~lpBŠ^�e9���V��!��,ql<dm���'�Z�*����[�(�p��[Ѭ5z��$�ָ�q����ԭ���命=� Xm�
;�Ts��P�O����L���ٿ_���m���r����Ã��a=���U�j*b���r'Ȋ��W��瞞D{!�K:�M��0�,��'ZNM����Xm�B��B���(�R�p��T~n��r��ݩ��MqN%�,z��W�=K����I@�a,��Jy����F��`Z�{Y�q���S@�x fe�l ��	M�|Qǈ�b�:��ǒ̉=�}G|6Ͼ����b8td�����:䭏���{LC��$�]�vJ��l�	�Z��G��#B[���hd!�X�/
&�.�Eyl�ys
6$P!B�8I� 14�`�
5n��C�����/)}
��8\�yq�Gb%�����0=��S?_�r/�����`�(�ݩ�Z��)>�̵QKXˏ̕;N���(f��`���Q��6�O�Zl�'�=[t��^�4yܺV+�+��*�NQɫ���=ՠ~�hQl>���\��K%Dc�ck<Y\M���TdZ����%l;��Uui�wa�t�NTQ�]�RH?^��?J#Ju$�ja�)	�ǽ���6g�e�*�p�Iw� ��1c���y#�mf�k�������KzS�y�ʄ1����ڞ	^��ز1��������r~&܎7��t���Yf^{Vct>�����
Ç{���y��5�D7��w�x&ë�!���{�e��볍���m�H�=�U�- �����Jܕ5�5ݳ�ԙ٤�(��KD���Q�Z�Ha�H�y%u4emVS5"��4�Q�[��̓|s'�<�}�F ��C����s4VJZ�,2H_nZ7�l$z��u�5E�-�ϻ���1���Lq0������L���s��BO��*쌑;Z$@G�:Bgv!ƴ7��xu3m�����<���,� n5��-Wx۰��gx�1=hh
�����:X�І�/:r���A4�]�W{.��%6!�j�
*�B׃5Z~v����}�R� ��0���Z:�Of�{L_�GV�%���YskMl�r�#�t�A���n�ё�P�q��Sۗ��T�J��d�p�P�f���psG�i�:����/rR-�O0�����$	{,2�x)U��X �kn]1Hz�r�eM���=�٨6ɌiKL���&�Y�Dvem)�di�dP;�z_�PQ^�-�=�hg�O����I��Y�o B�ܲ���
��(�" ��m�^Npy!X+=���1�����R,�6 �&��'$�;3^@;�Ŗ���*,O�t��r�.��k0��lxt�d�ZX�0&"��Q>��F��'d�}����2k����Ȯ[g��}��IÁ>{z4�sk_�.�� Z�Z?B����2X
N�� ��-6���P�K�'[�Ϲt&e%.^9�������$��GGR�� YX��1�:~�S��d뱰��#��,X��ƻ����,�Epd,�jE�E��X���K5�*Q�Y