XlxV64EB    7362    11f0��s�Z�?�z'���%�D�ꜷ��}������I�ZI\���rߪ6�QHV����~�9�l�#��<���� B�v]�X���T%�].nFD���C\�6�e$ɿ8a�b���ÿ�1�Nw�9���y�f�K�2��Y �!��酀�9~�����k<ó�%T�<Z'�[�ov������R$�s�t�˼�z��z��,��!�B�4���Z_�W���+��tz�����YE�孡k\�Ę�O{fz����8j����Tt��,mt���n����=�b���¼�]0+�ܧs�zu<�
�ږ�2E�}�`5)�xM
������tC�?� iׅ���� ?_�Tw?3��4��-��o� ���f�×i��Y7���kN�#�.?�sL��zq(�X;s��X�'%��|�$8��t�������hQsI�LY~�lX�U:���1�dWA*� 9k�ĸS��k�6Z���.j���>�a��ē9r���u��o��&A���v4.�����(���s9��s 2�bV	��s�Ȏ[F̪+�yʅ���ޖ�V��)#gͮC�\ �q?�fz5�r�?�WGj;.i�V'l}9	8�!�2^~Q֓���HDW䘐�ߺ?�-w�����ę�0/��B��3�/P}u��۝���;jn\��3cK���`��מ~e'� \rA�f��Sv�#ؤ�L��A����U��׾s���ٚ�ym�L��]o剿�{��|���-�Wg���B�L_ve��	�U xm�̮��X��x2�h��ǧ�6�t8����RiR��[f��	O#�o,k��H�8p���'\v^�S󘓬����#�)a35>���~��')�
W� y�-+��S���ZD$5�*{�_]k}���F�9�����[���?��|M۳�6X����Y���{o�JMWH,[c�v� &�s�U�r����Y�n�#�?S3�?[�]��ꐠ��87�p0���q~{YT͇Q��Ґ{.c��XN�4�`VY6��P3H�s�U��-e��_S��O��k<�~Q69
���`�M5܍��P�g�磆.O13V�2�&��Ĺ,�Ϡi�k�+4��g��'¡�!��p��;wz�yR�}?��6�N��4�CtR;�T�18��р�4����|g&��=���Y��S7��;��_�l�{�]	ef-�G�|2�p�wLOPu�'�4��)T�@,L����Oc�<���5.P)���^�t���gP�b��_��O�aG(�{ظ�����@lZ��1�n,�6v�~5R������KҘ���M9�,���=M�R�/_����O�v�R�UFkܙ�ñqM�_�S��6�T	��,���ȁ趻�˴��s��ﶎ��
�W��H�߳$t�b� ���)?��{�vZ�.X|�鉫R�uW��,�Dnu�J({�������W3]��R�H�z��5��O��f�(��@������-#F� *�Y'.y�&����Bh)�O�Ȕ"'JY����,�tmV$���� +ͭ�X?�Rq�<����P�r?�E�|��xyR+�_yWR�� 	t�uY�#��/-���+[k��h[V#���+�p���-}�P��`r����h	H �� |�Ax��'�6Q�3k�X
��5h��s��9�`��Q�cX�1�Rsŵq�����KS�냾Oem��;P�{�� �>�<�HT�`[�:"'���4��y��ҕ�Q3|e'Q��{��� +�c<�WU��q�m]�u4"�u�~X�i�-�ZČ2�n$�����:�v?�|P�����݇zIR�NIj�7���ƻ�-��.�;Y���'�3��ͯ1P�J�0uv����}x�\Ɉ,\d�q�7�%O�+�s�I����7k[�P�,D)��h�Qt�=��ei����,���˽�W����cp%�(+���W���Y��.{ݞ�7�t���^��@~K(�n��d��f�b E$rW�!3Ѿ��v�%�Oۈ���SO��-���R]�7��NsFt���a��ʫ��g�a��V�L�|�V�S�Q�y�O����Xq�^��=�
�9~��߰�[n�u�Ar5m�N���X0�e�eW�IC:�80��Y� K���^/f���R����R:x����ák?-�QL�̾l��_�o�������QH��ZR����=�#{gȝ�jJ��f�q�(�
�IҮ�z::� L����6!(Ǝ�	4Gt�I+w����;�TL9e�j5��Pp�k����j�H�x|S���ˢ6MtCBؒ��;b
�1��D���d�$D�=B�V�Xʀ��О��P�����@D��o�g2�2�"Q
I���Sj9��2����ֽ9��K4�N��� ,{O��I��|�˚`�Զ���v�735\L�:d%o&�	q�����^���.����R�k�C��I~㑼�x[x�Íggt�l����?���w#�q��֍�^|�h��0�߈�d��x�&u��J����Y����*��s���}j�~���E���zG��~�"T��u1���eJ�?���]lU�ȝ����o����j�!U���C� ��[�,�#u�� �z��}gu�;�Y��f�&��PM�4��G��Vӕ1~fpB��I�<����dR���"���\<�Օ�8s��T{�'I�F��?SΧ�P�	�Ɋ�q�����)M� �#Z���-���/�%]�#�㡣��R�����=��UW�@ӇDɞņ�z=�J�����F	ʤf.��]����ǁ��q�(xyWk�Lz�.�L���Oڟ��]��:�)*��Y�<�M��4�s��gs����R����霢,�J���,�Y���c�k	��p�#Ɵ�;������  �l2��(���Y��aw/2��+M1~��v�B*��i��@v��iH� i���xaW� �F�f�&n.W�ݚ��K6��wt��Q��+�RD�ʃ���y� <s��[&�5& ��f�K5}/>��]��`�j#�E���"�cq����[D���Op�*��4���HH��=�@m�LQo�>�V-VH�k��f����Tp�M�s}v�j@i�����hw�;Lo��m��{�J���ѓĀxzH�٘�`M���"y�.!��H�JE`Fجҵ�0Ny!���W��Yh�C��z#���6��:;*��K��5��c��b�-bBL���0m��}��z��2'*Aߝ��̹q��wR�Tw�s�����c>&}�g�0�­�O��oy�>1�LxA�F���S��C)w(t{�q�pmZC�v�H03��{���+��|��fN��WD��Trz��AJg�p��U!��D{҆�-Q���&��2��v�YA�WI�`_�m�x�m�!�c��k��N!"�o1]��|U�z�n��5�<� '��C+�+�V=Jq�A�%}����nu���} _�� �)q����y�U����=��?m��GO
��t*@R�+�fY��(�
�Iap>/�Y#��A�t�3���V��~�p�=�b�����}���t{`! ��i_�8
�y�o5�G$��[�v�2��ZC���� &������Y��s⏖sï���64	B�'����.K�?YCL;���+��k.yS�Z�#6����SqDGPl�J1�fꧭ���91p�e\���������\���0ύNqG��alz�O���Qt&�"��Uѵ�Q��?�pgH���h�Jc�mm��e�n�&gy�M�ׯ9M�-� �ڱ�ge�$��CNV��E�ڤ��e�$�#[Ӽ)g�<�����T>��W�=�I6UPl����JK(@�ay�py��Q� ��6w-�s����Ͳ[�Rw}y�C"!�4e�%%-s[�\ƍ%�����%"�Jy7�{i�X�P#��pq^~0v�ш��Ѽ���
��ĝ�@�svG@���h��a
�غC��l˕��:�pA��TQ�1T�S��_�t0/�9���I#��s[�M�5wtx��P��R����e:F��	of���I*��d���L�w��Ԡ<OY�����>"P(�ɍLw� %uU���0>��9$�⦩�W��|-~`��q`J^.�҈��l��X�D���;V�M��TL��(���k5p���3�!�x��W�C&�Ӯt1�����@
�z|岧���G�L���i����~���INv��aq�_Kl.��n��H��Vt��s	3�̯[��ȁeN\�����@w����)V(�NҁL��A�a�3������[����!)P֦ˈ.��l���y�	E��Zo�{Ѻ^7=�!"IgՊ^�mQD�d~�#�wJV��^	��C;�N\;�̯U���֬�(ՊWp���U�W�>�5L���+4�8�%b�__>ۆ�r.���YAM4�p���x��c%����F����&�]�3f�PC�x��Հ��
�f���o��Vb��N�e�.��]î����