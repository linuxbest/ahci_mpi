XlxV64EB    fa00    2f00i���yK����!���u���s�Y�sXE����1���3�X6�C`,��Q���0�n��I��P���:5�����:r��v�luV
�Y�8&{W��8Cr#�$�����rG_����D�!��,�	��*�Nz�G��j��޺��!��z��n����h��oJ���gf�#�L
T:p���w��QWN�e;�ܖA�O�#�ݷW�4+u����	4�g��I�~k#��)\�J��cV��>b�$�eOѯ\���]k���5��4�k��a{�Ҭ�ʛ��.d��BkC�.�G��|v�
|�Yz����ҭ}MYVc�^�;�?{�b�R.i�Ǯu ��S貉�m�YC�s�n�*�ʕP|��tP���kh4� ��}��:Gy�է�����P1�5d~r���>�p�dezu������������N�R7�����E�	��t ��ҡ'�tY��M�?+�{N::���f�n��Ϗ�o0�Y��9�JB���B3@Kڠ�Λ�S?!��U3B��H0��� ��`�!z	b%|�aCзt���#�2���$�:�7J!����������Z�8���H�S в����ʁն��}��޹��|����x0NH������h�WB&�⥶5�"�(���*�|�/@=��U��}?���Ь�� ��i4JXUc�f�����Χ�w,"�J/�Y8	�c�:���?��La�Y��m�V��4��AA��;-o`���gG����b�?L 6N-���.^�Gxy�F����`��y(��' ���Dp޵'���l��x��x���;m�1ù��iʣwe
6����'hW=�Md�� ��v�Bc��]P�s9�)�/�o��r)��˂�Z���7"ಈI=�y�K�
�PCi�$�g)�W�e��_Sٱ\�yO�&�Wk�d �D���(v�c�Ģ',�qP�%QZo����й�[ǚw����l���E#�R�lE<X��K�r(&���l���xE��͸~�ᤑ�@��.�\�A��^�`hޣ2������������#:!WNH{К����ES	�k���T�$������ґ��a�����Y�?R�Cz���>�<(��G�V�����4�xw�M�uI;T;��g��R`�Y]��k�`���~�ker�pmJi�:�t��l$7�9���
<=[���98�ّ�%u��^GjP%5�j�=Jf��"�����#&�Y��:�6V�����Z�,�O���ט� ��M�K���K�O����@�$���m���Ԁ	Bz�9�� rk��s�')va���C����s�I�j�{��:"y�޼��ق�Y˹����/���tG���ܸ�mJh&��S+�F�>�hO�F��[�2�ZIfp�ڑ��� �S�믕�:��;M��.�D�¤��.
����)B=u+�H8�]��Cߒq?{�ˊ>H��|��<,��P1g����/��5�Cf�	�,�y�ӥ%��1�_��u�E�����78�m? �P�WS|����<{P!Z|T������524@>P�WĻ!}��` ���	���S���;�Q�Aq��|2Ǐb��(7��B�!�/ Gj�WD�?��En(ߣ�^���q,��Z��K	�C1�R�7�� ���÷Mw�u4�J��sA9���+�.��H�Tb���˖�pi� =���С�G$�b-�T �i��r>�^]A� :n�,,��ޤ��U�1ɩ-?x*�jt�!��܇�gr��z3ɦ�+����H2}��r7e�{�5�����'FKK�:X��@�͵����=�垂)?��vVr��[/�{"�_vЧ~HL���G܈�2�`��5��`�S�.F�����<k�s�ѣ\�Ssοa3� \����
�EJ��ʑI� D"đ���Qcq D��K7(�h�9�ɟ��O����3]юᯊr8P���>s��m����r/!��ݟI����߾.i�Ӎ��B(�L�	��KixN���k�R_hRk�Gj@���K���W�zm�@��)3G%K�}`��Bڕa���Eo!��-��/�b�-�A�M��2��q�<'�/7�-S����T*�ď�5d�!�V�0��;��b�6��}��/��QH�	b�L�O����<"�ܤx���9I�5
!~�S��9̗�*�UF�/���8�6}���}�� ��2�jw?N�"�1j0��
D��C>��˗�W�#����!��`r%��:z�ć�F��F��ia��Hwa6�R� v��y�2�F	9�ԉx���"w�Y����E��bt��NAVָ�fX�M��]R��r�o�"����7��:�A�+�u+f�C�֗�])�=`���Qk��7�sv�w(��F�Txd<$_��'дQ�x�Y4��]R���͔rs|�$?`TfOճ��:?0x��ߋ�id 9��`G&��h8f�,�c7T1(6@R��Â|�!�C��!Tw�9w:-1�a�JM|3�B��޿�XDJ:Y�3\�� ��ƀ�N�(I跤0H��牊�4d�>H�֞��'B���޺9�8����W�4�����NJZ��"�:��_Ȗ��|^3(��J��zE� �\��5��äkP"-�K�.JȻ���5�C���Ʉ�,�0m�D��`'�Y-&^u~S��XH�"$Ϣ�G.n����.�ǐ�z�5��6�4q�����(~*��p?S����C_)�l����k�� I�*��ډ^EbB^+����]{dA�ڛ"�x|,I�^XGw�tU�c nQ�M>&��{H��`|��FG4I��b�ѾͲ�|�/�ގ&�><;���҅o\H�Y�b��҂�gׁ�%쬈�f���0�X5e�߽͘�:,C_k��{9܋�l��h:
�cz����.�z��ݢW-&?x������i�bY���eC�zZ<��``�׌Y���'��>Doj��C]�:���9I�R�3�P�W���qo������(������_J��S9��6�0ϴ]˅���Z6���mi�U�G�=P�IӬ_�N&fk9� �Z�@��c]gi�'��Ƞ�❝L8�n<t��^� ����Ys\� ���	���yW��g�-�h��Ns�R�[�vDJO����uT��o��p}�0o)}�!�'��R��A���6�nT{8D�g�3��_��reg�+����Ĕ�ɽ=�y��*���������<���cZChC�*a)wb��k�,��f>��M��0������ x`��~�f	�/���C��S$�;$������G�����<����s�଱a8�W� �vR.)|�C��A�W���j�bC�Ǉ� Z�zv%	jlᕗ�0p%�����U#�}P
`�=H����>�����z����m"IQ:���N��1_�t��0�v����"���s��ol�зRo/�_�uF���腜��s�WQ.V��������]3���2=��O{د���� �2˵�{F ��*�iu�"�>�gv���I��G���۳��s�cl�-b�0��p���pK9b/Qh�&����`�mJ&M��.i/7��S�	]��i���g�z��+p5UYF�`a���ًm���,J����.�'�T-�'�$pq�F�S
q?�����������|���|�,��:�R���'5Խ�����#T~��W�����EAe-�����58h��J���A���O��WV��r�N�p��}�_�Y�p�ò��z�^ӄՍ�USy3�	}�/�b��)���)���Ζ����P�)��9	�|O��ԏ��dDl�mU4����ɱ��]��6] �_1�=l�>I��W��o�!nt�Gz��a獴ԏ���u���桰ە5�먎���y�%<4�	4&��7����C0�z��Rƶ\ ���8RjLcA���b���t�|���:<X��z\*���HE`/���@ڵ�h���p"MJ����c�Fj���;2�+w�!Z#z�����ﱼ;uV8Oy68��S�z����?��8���F�yb��̊�������:�
�3(Qh���C5]4_TО��|� ���,�x2y	Uquڒ� y�~{DfĶ'1lE~�IM�8�D;V��jܸ!���c��*�� �|�V�$��1�MQȡ�Y��ܓ�2$ y��c#���8�ņD��/S]9��s���(������_�������&�i�=��>w�>q@��-'�99�+`���;�����!;�K[a����yī�[2�Ē0�"-ۜ,���#�|&�5��݇
%�DJ`>�X&�P;*
�-��3�4.����S�C��-K�g˟v��cR��/�e��8k�%�fs�C�B?��U!��y��~}�W�2�a������|��p�⧸��<\Y=]	l_٫�lS彘��֜�J?�eABWf%0˳'���Т����b�uՑmKq_�^F�{l��X�|7�tA`	!Ϻ��e4A��i�oit��:���=�)U<�>�J��k�wM��x�/�a����}�$�x��ܾ��li�"pHa��(Oib�~%��ϜAKGV���D�u�=J!���R4��M5���]*0��?�U%�a��(�ۑ�|<���K�<�?�c�<#���X�X�'�&@8*���4�o���C��є+{W&�6��C;�ȗ�wu�<��C��䵊�� D�xcY���Oט;+�\�
�`u��T�}�ή�� 믊�)L
ox��j������F
����cϧ�9���58���)c��d]�&�1�dpB����N}#���y���r�ºg�dR������̀��/8�%f[�g�;��ͯ�������S�;,B`�d99��Q���i��Y�m�&�0�),5Z{*y����:z���/�k�w_�������)����`9�'��v{%ض�P�3M�Z9��Լ��o��uj���a�v�ϴ�=��-��{,�����F���{�F�#����	�(�:E�W}��U|�b�	Y����<�����<[�g�`"����h������-����������!�L�,#�n��eU+����H�Ҩ�Q_���;�H;�J}1I�� �`^����y�otO<+Dڰ\sT�٢��
��>�W�JZh.�T���o˼*��`��U�٘��,V
�Ow�	$��j�Q�����4��@��M|X/�~c��ۘ\L�}���%��Zo �-�o����,�f�j�4�����7������f\'�����4VqFa��>��8Y��Q�����b��a^=�UY[�?8�:�T�ƕ]D<�|�'I�:ŝ���3���A�Vpd��9�:v��^���p%���������4V�V@RirV�ݨe߄䳟5ӭ�F�.M�"��[1���W36�[�'+�H�����*��U�i}�Y���Y.J�d�Q�ϚGX�_��\7Sc�ߪf������f���݋�L����8u�����op'����D�F��ǶH$��A�l�����{�9�#6�=0����K�����K6.�AUf�r��K{�E�	�X�ŭ3.�aMH�¾�-]P���`N��<B�5�<);���:aLw����R8�MY������T��=���|D2���b��ޖ�buV�|=��u��1d�/6��}3#�¦M_>(e��/����c���Vc*��kE�HJKV�����yT�4U�1�����f��P>�Մ�#��j��0�ޒIA[�Y<�B[���sYD�%?s�k�2)�Φ��p�@"��œ�Yn�kZ��x*��L�
8&��ВC�����ʪ
��-]7X���
Ģ����	����;�|c�<�]P�-��y�3?O�$yg�?|�)m�F�In���dȅ9D*7�����5���/=""`�%E!���w��m�"@�	|bK�̀�  ��N�oۅI���p'EUͅC3�E|��]�Iz]͌���a�	�Bl��l|>1�w�&�k@����l	X��dю���q�R�Ud�@�У�!Cn��W�`
>LW�-�,�3{���4�k�Z?�
��o�\:>HY4Iz�1�	C--t�IN1��xY����J&�CB�h�,�\�^ce�A��pډ�9Z��l_bȃ�%W�7��'��`Mϕ����qe��v����"��ll�L_0J˨�;�1)l��~�$sᯚ7�B����������&��r�� 8��շ�ۯ����� r�'��)��չ��N��������2]V�mo��C�C1+6��v�(�_-:j�Ԙ
}��d�Cuo_��L��=О8Dg��R�]z(33{�+Z��Չ��16#���HM�v�뫳s�ˣe�`�"�"���M=���k��m����I �}�Ķ]q�jN��(ee����)��j�~�Q��]��%��񿖔�i�$��^˫4��U9@�t� �|6�#Ҭ�`�43���	��K�Ӛ_��'8Oa�ۜL�����pX$qڦ�����1S��fe�>���^;y��7ͪ���e6g�J������ťvל3��JȬ!gLȫX٦
�Ù��q1�M뼔.\��&r�UM�S�0X�\P�We�yn��
Gg���Z� D�W�mG��3p|ռ��U�[9�����Raѭ$p���W����|�p���i�"�"a'kȥ��r�m�\M։����M48�%�����c�&�쵧h�}�(m��2⾐�d�+,�t�W��1 ��]T���s����J�UZ���A럺NC3�*�5� �jE1?���d 7W�D-����.V����w�Ï-&��^�_�{�+�V�y��`p����Zf�D�1�@��\��,��q?y�T�W��]��T�ow䩄���� o�'��돮��(�� ���#��+�Z���l�7b�j��l-�p;�.@��>� j�+0Mپ޼X��5_q6�(2�k��-[�hK�5����=�r�:N7/^o6�<6@�n����>E���M�{Y�ς9��d{cI޻�>�~��5�w��\ω�p	���+V9��1��(к�5LP��9����:`
[C� ���R��g>�6���V�/��, ��l��.��Yx�����X���A��e<<+��bA��u�Q�&D1��:�/��7�{ܛB��2�`HǧSP���Qz`��H�
}z�mK�A��?j�%�_ݪ��N��e
��y��~�L�돣��(��="���h�3a߼Ԙ�M���	kk%3�� %����]$�~;.���|��["5k�J츭OY�[?B#���[jP=!|P�n*� ؉q����BMz�Q9~�s�)���|M�0Llf�@д�f���`"�'s��"0�]b%�lq�d_~���V~s��W�u4��s��+X����6ųL�+ٱG8X�:%���i���jr���;��"�"��fn �	��Ñ���Gu�U\y�T*��<ӡ_�g*l�سeU+6a�WM&5�pͥQ�*+����ܢ�)�"qr`�s������*�P�h�$�Ԭ������
�^� ��wZ�B���=c>QK���}�������"-�=4����\錎pxC���P�_v�,����F�;6��f���||�82�U�{�S͇�����O1����)�A��a6j�����3��w:�';߃Ò��R�K��b�N�0��� �A��n�p�o�te�G�J� �W.ē�Z��'��Q/�.�fǄ���
]c���e^"��J�_C����PRJ
���F��|�`������,����H�[v���xr)@�Y��<��A^�i�|N>������BK����B�ӄ[p�
� K����f\n��x��h^�Y!d�S-� �h{Rt���	��������#tL���b�D�T�!#���	�0�be���ul��tW;�d����Y��x�خ��}ܧ���rʃ��n1�>hC"���F!QţeU�2��cgY�9��^9���3E�&	P��Ⱥx/��j��MYt�ww�:T)Dƕ*b5�v��҉���̳��?](��7I/qD\��@��1�nD!��e�L�ݜq@��J�9�[jl)��M����#�B6Kx������������F�2��P��;�륹]��c�Er�1$ �/�b���9�*�������iG�S%�<~�'��b���79S��P,���:����匐:����!�T|�n��m=��%����6�)֥�:!ۜIL�3���T-�#52-o��ɀd�;��/Br|�M,���fJ_���S����-?V����`z�"E����"�?�{�
�?�M���B�D~��:��|g�ɃlBa���3�a�\ܵMZ����)&���<
R�f��K�(_�b�_���coat�|�
�)���R4�^�I��柅$�L�9�9s��"�nf��t���IߡM&��/:��	cS�0j���͋�m�G}^�^[_����[�M������&��>�{|�����{�z�����t�	F�qd˹���d��m9��Ƞ��b��#�v�5�4�	���~��ZV�^�t����{M҈3+�u~���P������b\�y�񇤦� L��'�J?��`�btA&���Ц�$��ޖ��cU����"�s��^�Z�p�p����4 ��Z���A��2���q��=4�տ����$p��������R����=0V�B���N�8<S��W\���p܁�l�8d����Þ�w�жQl_RȎ�N� E�<^k��T�샚a�_��i	3Em4C��u=��):[�$&�v�9����<���;̂���I�B��?�L�#E�|\yq�B��丷�?���no�Wh���5�s}����k��MR��Op�nyF �:��$¼F��%�HZ���d�E�zEz#�Tg�f��6/��rf�)"c�Z"������x.�ڊ�,oe6[��,́��Ӭ��h>{�D_��"�$ ��Fg��(�&�����'�ԋ>��ܠb��u7�5Fh�+yeė�c;�|6�Q��a+�?iج���Sv ����@g�P�}��UU�#��Ҵ��^_�-X
QoXw�Gt�9Z��S\7����$uSQ�L�g�ͦl�*��3�t)��<�,������I�q���%<�>=��GT,��خ�K�(\^�V8y�̵(�r�q��X����B�ux�5���/e\z��y@���%>�kB	�l7W�+��8�!�:�(�.��4X0N��|�*7X\�����/sh`����QwI�M���y[[��$������_m_o��Y�x�K?�����Җ}J�0�OJИ���0�Nj��� )����D���HI��n�/��|Y ������͎a�ޭN-�5���5t�[�ɉ�s�*��Hsx���/=��M�^��ߛWU�����!�� ;~t����������JD��a�~��
ՔF!�'��bJ��3����n�ʦ��ƽ�ԓ�[c��s�HKR��7��ܢ������b�v�q&b�dv��F���<��p�ǩ��p��Jv��+Ƨ~NHJ��4i���.���K.������63���@?�K�j���#�K�Nϼ�)��9��]�Ք��䈔Y�9�.�r�_���B&Uи�a���.�G%�j��<�� $�8Qh�8��{��y(��(Q�/��>~lĿ�D$7���V��(���W>A�/�h1�]|�8k�)-D�d�Lf��_ބ\� L���}�e_$��a�����.��:FX�xC�3o��(�/[��o�&�4!�C3D�����nGJr��O�覜��f��:��NQKX��G��}�s��}k���r�1��\E�¸[�u��e���}Gh��� ��u:�<iU�����}��	��d_/x���h$�R:��o�uYi��Djܖ���gYk�@�˿"G���)�N�>$�B�����v�[nR�m%�N�#V���=Ϙ�����Q���_l�-҅|ONK"rii��ϲ�@�qO������5U�Q��
��[;r�Ho?���i��� a`s��Z��H%�nYygM��e��I U�oiJ�55V��a�1I:�`�T�Bqw(�@J�uհb�+�)���
��y�Ws�W�)�3Ob���
~@��k���)hbX��YK�yZ�
��4UV��w��a�<��߳pτ�׽���EEEB,�tK�һK�y�iZ��L��z� ^5e���6[�I?Ӹ�@���@�{x%P�e�@��^����mi�Cf ���M�n7��	���i���C�D�/��6�%V;���4�{���N%�}5L.�H0��G*"JY����}��'k�qKPmH?���!F[+�%s�W�C�e�e�p\���iV_ 2K:N��G
/!m���yҜ� 4�@�z�Z��«�:$]���#�0&���-�Q
6��CϪ�r�O�8_�,�BBsv��m lЮ�%B�����z⭹'�W�I���CE��G3��BM*��@C����B�|"D�*�^�f�^�����_S�;��e��L��\�
�b;ߠ4�,�h䞰М��3e�@���Y5���n����2 �~Gi^�Q�(�@� �6s�V�8�?�Hq�5��%���a�������"��nk��dx^�Y[��Ά�ֶ��~%��V����l��RF��U�~�ݓ���i�*���6#3��{I'#;G����I�m[�.�r��?/��?�`�@��J�s� ��Z������1��ۗη$bJ{	)�\��3`g����hs%��Z���Y����<��ہQ�:����e3��jT�!�K$����X��u����z��	�C���3.�Ƥ���zV�ޜ7V5�r�Y���~�P����x�W��;�B����0���)#����0�p��}��zۥ�9�0�G(.̎=�������|����� NU+F�Sp#�r�L���o0`������*�*�1Mp�-���J+M�lX}��9��y�'�j��������˨(Un`�6�D��W��z��/<*�������J�p����*��w��X��ڳ�W�K畒���\b��4aS;Q��Iw�O��.��_�qQvQǫ�Ƃ�C��2������	~Vmy�����9����}=�'5�\�e�0�� 3?�n��H����6��/�<�o}y�0@0�r/~�v���ܣL�i8�����;o����\˿��r[��x��<û<�lyȈ=�I��jz�5�5�!y�TO�@�O���5=��F�qgZ
*ػ�:^Ԑ�o��3)\�y-m#�0����. Q�K���Ѳt�r��&��0&OPS&_r,E�B 6~�o�_ן��.��]�I�j��c������-؈���?F;��l��sNĭ�SF����E=��F�����}��rˇ"�D�5^���i��֥�ٱ��8b��%S�S4\X�g����T���4�����N$�5�˛���74�q+�n����,�(b7(�P���.�^��y�[�� t��3�y��xNw�!N)�\L��c��e���6ը_���v�H������wtp�]t���f��r�v�|�(�0��<�!�zm��tBu�8{�n�
D}��w�C1���6'%�����} V�{F���� ^c��QuG �fo'b�[]8�����)�W͘�J͜�,x�O��WՎ
d�$3eNh'EU�ǐI5>��ԩaq�B�t���Q�~����4��`���L=,VV��qV7�=Oy���������Q�L�>�NdZ
��?an�1��S�Uż��<��H(+��κYYOD0XlxV64EB    c312    1fd0�_E]դ%t�+G�Q2R��}_�LH�']����"mSN2\���\��sj ����J(�Hh�)��J�G���k�ݒ��x�H�5�n��,�SeX`��G��+G�}r��zW�8��(:3±�F�kX)׽�d��2��.�g_�mu�4Ԉ2VQ=Y�S������������`�-T�`HÍ<&S6ʑ�բ�s�����̸� K*�rۄW�uͻ�6�gŐ#��k�reZ��-&]�gD��G;Dno���v�0R�`��PV�����jfh��SDc�Ix��U�%JN WXr�
�O��-rL���;̝Vk�����Ӈa���n�8��/�S �)��]�鯲
������F4-t�6��{L�_��Ip��G��A/��gY��$e��G��d0��&�_Nbh�x^bw4R�"
��[u��/-�Ƭ�%U΁%�#`���dA�ǹu�������r�ϒl�"�.O��f�5��>��m�^��� ��QUX��f�!�X_ɍ�+lb�>S��m���5yږg�t��
ô��0C$D	KR�5mP� �Z��ɯ��H��P&�s�a����mK^��߯L��u���+��ED6�Ԏ>,<����*
Y����7��&I�5�6Ur�0xlG�n ���ɀ�n�=z�h-8ZPw��r�a�Q
ߑ����ġ����4By��hIHM#��"�T���5{�%��7a|�(��p�*��gǮ� ��<+^�@���\1�ut��sT5�� ��ӹ𝰙V�pq�#�Ԣw'm�hu}�G�YN�eӳ�_8���o:��$j�F	Ș& �>�{�;S�: ��3&���#n�y����B�����bK� �{	�E���ݲ3�$~���E� ��o\�����h�n���l%B+$e4�U�k+& 2�u���K�yLS�Ԫk�"o(�>�ξ��)'�#�=�lTi5
���zL�o���g_SOs��vF��\z B���R���e �:�y>�a���8�x�[�O����MϻYlN{v���߲Ia�i���~"�*fV`��9�u�&�/_����z�i_�h��Xl5����̴2�M����q�*���8"Eg�������-ҲY�, ")=U����j��\������/b"���9���r�X_b��H+��x���/�B����~��?��,Ky�Z:KE+�dS��y��{�{ڴ�m��W�㴫����m���&c�m5�O-g{Ϯ�^��,�w$w�O�]�#�( .��M(vw��t|�{ުT$�}�x�8�ق�.�6��b6�/�F_�:SLP�W,U6�Ƅ���s�Q&�6n9�%>a�p^�vG#|��ot��O��C�.q�3�V����� �����S0H�ݗ��>޻W�wz�so����%�D�d� ��������a��" �9�D�}�Q/��8���N�f�ۓ���<���H���°k���}�β'w5v�z����-�4�٠�Azm���>(Gr�r��A��l�e
8����R�z#2��n�,|��]�b|z����5�_fI�I��v��sƾ�k�Ykd ��1<�����4H�}���l$[Ut�mR0/�a�ξPr2�:BP�qˢ����x�F#6����,fm�?�@�d���Bq�ͅ'�l��(ߥ:)�m�$�� K� 6����.�ʠ8�w�_'���:c�`��Bh�o��!�:W�{���F��L�+�T�lSi� �|.�t��E����ӹ�#/�.�v
m�kbCqxKn�p>,\�c�S��jSB�dQR�ݼy6�����o<�r~=�@4Gsx����ɞX�-��~6jpL���ܧS�c���7��j�=��lM��w�	��i�Et��{M���DXp�y�v�p�}����A�%�T���}D"n|9�A*F�lP=�"X��V�#��"�2�M![��UP������y��$�C���ͻ����xi!1�;�Է��N�A���i֮
�^����~���TN��z����%Tq�5��!x$�X�3i^$�-[H��܅^VF�j���xc����p��r�WT�g=��CD|����嫁����4�I�%U����#���S��k���_-��_*s?�ea3�'��pL��1�*�_v�M�(]] o�&V��h�� (�+�H���x��:l)�,A�=�d�{fsj�L��)=ʱ����ů��O��Y<
�"D��A�E�:&���D�J����F�18�@^��ct=y�E*A�}k��[����\�<{qY�U��쳞R���N@�����0f�WY���R����%.�Ӧl�Q�IC!�E?Nϼ֠�/}<,u�����>L�i�����<$�VtE�DC�>I��N�ڼQ
���8b�a"p�k�a۹@����������.x��Վ,K����V���f�.{Vfr}��#i�T��@���2��b�hGI���|>n6����#�Y�Q�1ER(5=��	�(ZUE3D\9Ur�xqI�����0���>s5~�˴n���Q�$\]�����R>6{��z�C�K7����5$(W��`����y��O"��m��Kq|�uhp=�ɘ*��E={-e�/�	�oL�G��l�󈖓��e�$�������Ȝ{��l�񖴿+�Q�ۥ7�\3�T�,5� �f�x7���§�m?���x5S|��7)���`�y��qzS�	l-��á"SD+���\��?r���ԃ������#ERB����h�>F�я���դZ��N�A&љ�g6#��1�J���q;�ꚕ���B���U�s�~�� �����b�v�	�ɹ�kS[�h��>�����<��FC�d>I�?`+P'N�j��#��-@�>���x��~"�3�E���Kg���G���Z�Kh4�6��b��Z<�S�ҕU��U�_(�td����/8J����^��M��l�6�(=��J]F$qN7 ��I�����b4��' (F7VpQ)6rz7s<ܞ�c��ݙ�~��rIN��s��ш^U��p_�-��r٘�Œo���/�(�y1��:x�y3�C���GdKe/z�,j1�^�e T�E&�EVv�ꂉ�
����؀�#��[��K��owN����9J���nǁ��e��g��y^�'l�{��i"���.��+W���k55槵aO����|�L���b`����"��b����eG>cR+Q���q���A~��LA>&��$&�qHu@�Z��k�B� ��\@W����#s�B9:^�z�}A�f�S����s�l����s��[��_&g%�I�� ��<iD�����<.�s�g ��{���BY��_�9�� 43�����tV�9@{�c{�6�F�u�
�� aI7�4��Z�A��*�/�R�*�ݗ�sK����|�N��
胳@�^�����
m~�3�~]#����Ֆ���2u�pn&������1���!� �����/KX��G��Q��I�f������F��k�&sCǺ!���ж�!��(�@mڡ�X����|�6�m� U��n�?%�=?�Qp+�&jſZ8^�?5K�����oQ;h���$m���$�[��P6�@����2tl9����ﵓ�D��G�+[R���Z�w��|?g��|	��Oj�H4���ŀ�h��o���{@
�	z�~y�=�}�j*'c�X��,�[��ݰW��:�X�a�t������rU�qMM��ոͨ6a�z?Gi�1V
م-Q'ߑwVF<�����jŎ�!!�
t��A�(�+X��fEU
����8��(u�e�e�v��L�`n�~Q�rt��t�≲��e}\���3^J�8���H�(�[r�~�@02G$Z�Ш��u�2C�Tr�dǆ�H����I���:��g�*pZ&�b$#��7����7��J�8J wۙϘG:&�u��X�r�œ��� ���0%n��qBu�4c����Z�J#�p�&{�"�ɻ����!C��3oh��^�k���Y�g�!�a��}��U+a3z�"�p(����Fʃ!��Ge�6��y�Ϣ���� ���O�y��mn�"W�� �j8�&��VbM_<�$�\r�DhoN�2m�!@]��}��c���׃,qO�ZLS�|����H�Ҳo;N�B����Rl���*DY����{�@~���)�����XSd
JD���Z ���ϯD3~#8�E��CC�g�p\6��(��"/��R�2�L�M�̳����^��dl3�$�k\��:)`��D9z �jOny�KJ�9\��s��⣜�N�'�ׅRhJ�+�"�5�n���q��C�^3�r	/�o
f��P�	4mpukt$����3�yԽ#���l�d�˫�ؾf`��G��=�����\�^\�R�l a�W�#(J��A(e��8|)4��uU��;�:5+b������R�%V� oH1
��%�_K���tP!h�Q���q�>&ߔH��������E���l{�^#�3碲Bf��׈���FZ"(�úrJ�Nu��y�w�㼛��؏�[N%c��%n�l��Y|�9B=g-�0%�S��H� ���F�`Ѐ��2��e�ل��]���I75<ġz�����G#i!6H
�B�o����O���]M��J���W%�����"�#��T�qH:��߯S=��t��L?'H�,�b��,�[�mI���~����/G�4����n��x���ͩ�2�,�}Yf�y:���P�}���\��Ju#�i�3�-�G<];E�?;�����͡2a�@���<����:�!�S����F}�ij�	%!K/J[C$;LU9�3|hF6E�ܩ[%�O������i�(������B4��{����b�"��;��2RF���x>C&^sC����k���1�;�L��4n ��Ȝ���Ҏ�Te�9�H�=�����&�h�0��(���e�����Ț"'벜�.�G?��}=���Q9�6DT�ެ�|�<��0�Y���Ȑѡ�Q��V(��2y-p�?B�!��R��~1Z&�@3�c"����=�̙0��t��v=��}:�= �s�2L:����d�٬r���+�&6�&ϻ���xe^�>��п�P�t�!RC>��O {�K<9F�B����b\�ܰ]%<V������I���lqi��Y$��f&�U�K\Y�d��F�/�#���U�;K`�\��$-w�y�A��с��t�Sw�}��B�ԩ:�we��OL�T�@�q\���~*�~ˁs`�z��F��K���wU�?��'�`�K���و�"�b'kW�@�w��EqV��?��s�Z�)��{��n-�O��k&'۝ m"�e*����!8��H;a��$	"!xZ�0��s��ֈμCK!��˼�� ~�T�O�qxs���"#<_؝�	эE�Q@M��)Q�-�����P�VmZ^2�\�%����*ܒ�h�E�%���7��۵14�!�=����NF�R^�Oz;2�]�T����)%��"0s��'6y{�w����8��aVN�ˊ�Z�T��6y��Ҕ�*,R»K����M��x�s��\$�}�g�.ob�[V!�^E�P��Ӗ8���+�eO]��_G*X~t���}���h���ᴻ�&R���vx��EO�J3��v�[ "X)�GW'�O7Ĩ��љll]��j�`V�)��o�Yk�0���R(Q��UY���o��iܸ�Tv�����v�����,��	�Yr�ҳ^*�bS$V)�0H"iS)f��tbo�<x}������%�,y�3�HS�!�&��|�;��>��!�/��\��_؟y�+\�P��Npc$zi���������T�;T��X��#RN^�ۣ0��x/�O���"s�2z��9��0��Qy}�0`�a�^�|�����������'ݪ���<�0k���?lנ޴:��l� ��Qtu$�r� �JWG
 Ǳn���E ��%Z��6/��H�Ǖf⭯"�l��,��Z��$������Φ�)$���m/r���c�)w*�}U���<9A=mRX�����&�g�	�M["�'�1A���{=�%�Ɩ �8�j�C��*r|!��%C��e��!�ゾ���z�cx��F��\<G���n��%u��0�����OX������d��k*��`4�,�����#g�`��3Q���?��t�1�O,��sh��#Vɋ���a�� ��ć�&K�~�)�G�z}�G~���֨F�xK��KЈ'��ǒ�+AO��E��Z��k�]Lm`��K��΂��'��Zv���U3�Wj��_$�j�T�vV��Q��������9�Fz�k4�sB�uu�d��S�"*H�a�4v=�F{ �^���)���T):�K㬂�I��>�$4`��q�n�ۜ��$�]��NC��	,�`���eD1��z���"[��� ���6�>�HT��jZ��f��FB���V���|d�e���Zr�D�j�
iډAB�v��f�i�?0�Q���)
lb�	t'����G��.w%��z�G���;��;������^M�]3#'F���SXȴ� �!��*@��{XU`�~cq��p/�p��8������Ag��F��ٟK�j]��q�nk8��l�⣚�5���]0a,&�t�o���ԩ��_�c3y��ұ�,!�y�v�G'@\lʙ�T�[`�lv��
#�j�]<�;�\ը8P�l6�l�)L��6D���� �W>��	f��=���ϯ�Cn���v7��d��b�ݨ�w
<\]B�k�C,�'hOi�y�4 I�$�lm.�^��!���G{/-�u�$x�:Ew�ja���{�7��ڽb����w�O+���nuxY��D1nRC6���؟eg���V9/2m�dZ��WF81���<N{����ǡ��7�U���]�{^���
�"�j�t����Z
0a�`�O���9�P_�I�;Qi'̋�Ά�gn݈����a�sGggo��(#������c�MpU��N�(�O���M��=�`���+[�K�Ӓz4��(R\ax���˱����,�.��sͼN��+����C1��?h�Es-�^��h��`���j�c_Zb�p;ۺs���.������4�^!5�;Ir��2���!��7��[�;��;��J$�
kL�"B#:�	����ǁNU�o�����6\��e�B7?N 4���
�� �9R�p���|��M��������2�z�k5��8��L�8Ҳ����`�yH���2�{+o�G��w�^'����8����W\��w
�v�Zv����_���d�H.�љ���l�pnV���y7k�h���Q?h<����8�YG�?�{�{����%u�����e<1r�zQ��a:��ȯ�q��*�)vɉb60/ԄK#�l"t��]\&��Rƹjl❟"c,Jo���_%��R����(�I!
8�~�aNe��
A�c7���\�}&vϝ	���2�)�.A�g�1��O[Z�o��b�j�@������Ǘ����9��AΤ�g%!�������+F�����f�<`��-=�0�WƯ�/��Ա:�M^!Y�p6�S%�w����r�/8S��C�[������&�W
����'S�t�-4Tռ��=�	����q�C(m���8w/'&;�E��nO�;����F� �	#�w�r�
�l��H��xʉ鎴�s'�wN����&d�������-"�@L�,6׍L-k	��K��b���[r�:q	�k��%��HN��������A❊z�7�M���G�!C����O:��L3d���lfVs���4$o� ��Lfiw�-j���;:�*����7�r�R��j΁�_X]���P��H�-<9��,.�L��׹`6�qb�Բ-�J��
��؈�a�<[R@��x�G1���^'�l,uO/6�M�>��ލ�`����Ni_�ݔ�FR%)iI��e��0[u���u�1_���x���p�Z�O�кah�/?#�r�
p�^M�~9P�0���)�K��