XlxV64EB    32c9     d40@�e�m��=4%�ߵۻ��q��=�ws�`Y44"����"�=��(J�h�D\&�L!��n)%���օ/o�U�"q�Џ!D?�0���t���7A�C��9<����ˬ&��}��U����o���3�}Zz�f1_��Z���u�%)��p-�����\��~έ�;fp�Bm]v�je�A�Υ��&�"��0�!c�8����
�nL��ǒ�&��(��(��v�	M�|�e�8�ͱ����[�T��_L?)_+�ٌ�Xͫ��Q��G[�Cƛ���A�9�TDQ}�i�)�B��9١o)��|+��FBOd�p��o뙪���LY�G�d
��c$�k�Sӥ	�A͓�B�纮��jH���'��b\�
D��;d���{���	����� kڬ�]6��ɐ�.L����Z����by`�����ֶK��<�㽼���'Av�&�΍���}��Ǫ��K$�Z1^0�J�'|X���yji_��D��ʪh�J3	ޙ�ܓ@!`��lH>�o���7 �V@�J���[�Hi�2 ��������&{�v쨟׻�J�rA�3���܇u�^�K8-�)F	f I|8~�����'�S��4z��/i�a��tC����|M7�R��E�9��5���fK�6�������E�|��G�A���e;���U�ڨǪ���5��[0B*kv2� %�l�`Osi���T��喬g �x�m];ۋ�X�*�5�Z�I!L�偽��՛�������I��G�bF�i�T��ԕ�T���lA�͊1�;1N�������@c��Jk4?��+��Qvs̩�`����bjӲ�H{������R�<A#'&5R�j�CգC`���/�a�vYw�+
d�8'-o�:��w�����n���J>�X��Ъ��2š	���B8y�X�S(;pE:�� �ƽ�G���Cِ6���&�G��hes?]��#�AV����E�kW<��3 �Al�/������q|hј���5%)\��y��C�>��7�ᥢ�ý��)�����Z�P�-9u�iĀ?sT�C'M7t&M�o�\uҜ_��t���jK3w�-_��J�l�j}�9��A�|6$�>a�d���n�����������P�3�����&�J�O,�rV}�Ktw�C#<�+�m~�Z5� M��#���9�b��U�^eˆ���/�e3˷�p�vζ���G��L�L��܌���*OgԽ��>=�A��35*��G�������?v+�)��/�Ӧ���D�T���<�LJ(k����
&�3��ڮ�;[�Z���ч�E�|k�fu��7��k����w��W>Tj�G^#��f_�@��,XQ�_P��^���G���L�&��/�z2�{B��Mc)d���-�JK{4~����X�,	�~�ʱb��M�4Ǔ	λ�4p�5��߄`�H�vA�JZ�꼁���W��%%�MP�΃R�����Q���8��#�"�˱��_�"l��N��m�(v_�4�:c��Z��T��=��s3�&i'OM(Z�B�M%�(}1�ϵ�ތ�JX��5m,mr��֍֌l�pW������u 9o�w��"��9�߰è�;��Rbz�g��f��E�=�j|
2�i�R��6�W#��	pJ���2��������V�O��$0��}l��G�K��f"e�t��8��=7��b_XtJ4Yx�|�xѶ�w�@t�g~M����p�ǔ��"��N���ـ
|�@1	ݓ�zB����������ƽٛ]�W��ub�F�D�z�b43��q����H���j�U.�]X�=�e�����RhF}�MǺ����{��$��������&[�� Į�矊�wZ��tr����kt�
��]�׋J-��A,���GX8��`�}�t��ڕ��C4��k�ce�S�x���?�{d��bm�F:���mg�-T�	O�a�����P���zK��X�ES��_��	���пH��n�6�������<��ߜS����~�+M��D������*���71�f�����\��g�	�k������b�@���E�:M�,i����6�e�n��ŐP⒎ϫ������.��GW�
�A�rN��H3`�]0u-ˮ�#k�L�9n���\�6jԷ9�A��^��I�d�'V>��_؃Ml��!f*_�q��3���M�5��]^p��Tڮ����X��YSJ�?,�z՞Y��.�S����(g$<�R���cg58�Z<@��8�J���r�Ĭ����îL��.3Z=��4^�u��ڭy�ݛ��d�6�{��(���~�@��h#�~8��T�(����R�+�rg��J�<z��!@�0��N���#�ا�o���(Cc9��*[n��O����ϣ5���C�P��7������:h!���t�jӰ�g5���>ω"���*�81��ª䡼���'��ze*��N����]P��zf�aOE^�����{�h��:[�=��k�I"�`��A��5O�L�A��� '���a���2�9�E�A�S�C(^u�+����zΎ[U_��`(��QȚu�&����|��Tk��{�7�v����u{wɡ�B��cI�����	cG��U=�	0�U�7���j�zo�R�YlZZ4��$�DM��Q�U��Q�gv�Nk!�,���gFG�"����t�:~��G�VMD����\/�x$�[�<]�$��_��T%ǉ��2�����o�h>��]�+5�2ڦ����b$(��,���MJ4��iq
�}eE�m
�Z]���{�0�}�-�V�l{t��(�?�l�x����ΦJ)�LAʟ�<qÇx`�h��h(+�VV�)��B���H�#�E��+а��U_�۞�H���"1��ܪ��~��η���%�#��V���+��#a�ۊ��`�Y� �|
S��;�P{��Z��~wD�p
!��u͕R��V���m96�qqJ�����3��QBH!��T�M�qp[_)��eg�&�8i]$�����i�bL���g�ݷ���N񿀶�J��q�ZU/�*���s����&��SBK����'O\1:�����E�`.65�8�9o�Ԧ�Ì���§8� T�����DjǔGgl@�H���"Ɛ�;�����_
v7ק�l��e�x!3/9r�=�����Lc>l��mW����VK:�G0<{#���v0/�M"�|d �/�s��EK��I�W�z
=��-Nm�r =�+�����adQK���[e���R_�:����u�r��ҏP9�h�p��`���YÖ�
�l�p���{���E��F�