XlxV64EB    5295    1510H$зr���/�/��Uts;bp���d�m�\ྡྷ�o���F��P�r�@d�&#��
�1���v�e��@2����xQ/1��(U"|7C����ձ��<�QӃ$�U]�/��#@��r/ߏ���ƴHAvT���9�yt��w��dk�������/r�kQEt�|d7!��+��H6�1Z��qn�խ���{�������x��{v��n:T�.Hʛ��AxFuvU���&N����plYM����5T�QZ��М)�ǘg�M�n����.��n=R9�c jxT$WK^��%��t*A��1�M`�l�2�V�!۶ex�7��@=��!5x �1�L}Y�³7����,��n��	8�c6<�+E�0֏� !��@޲@x��J9?����{��f�g����BJ/����H;\�?�㰐V����$x��~�s����<k�2�߿}���=�l��y��Zۇ2��C�}�rj@`Qm�/)�~s�p��}�6͠;a�|��N$�N��?ɱX2G}~*���\�Ǟ�b��gNr�Qǰ�&�}��#�%����7p�g�.�s�_���s2�}�y���4B������%~]�Q�$In�����
m�����ѕ�S�?Pf������.x�s��u6�O-��a䇕�"x n�n�hi��sW\c���`�bf��d(;���
ݥԬp�<�~_��gE���A}�]�s��2�V:5}��Y�/�^�]�(/:�7��|�[J��p{ajyq���
R�O�~B��p�+�[b� ��k�j\q���U\?����8(1E�#d���m����!�p[\ �3�O��d����m�Q�4��;�o1H�Iw�m��;I �)�c�NZ�����Ő�/i���O�	Ub���_G#-?Ţ{옥���/\+=
7�Cܻ���<��F�ٟg&"ے���r�'�sQ�u34�d#��BC�.C���{�9�Dmu�2��X��~�L}���_]���}��x��!�F���©���=N����{dEWz`��^T$g.�q�]���0�G��l���'��k�9Rx�]�vo"����Y`�#�Dt}o��`��/w�����U>�0-���ٟ����L^>	�c�@	t�=<s6\<���@Оep�*�C��/d8��KQ�O��`i�4ʳ]��!W'���M�0Pj�����;�3Y:ǅ:��Ș�w���t�\��vd�Y��cջ3m��T.N��v���7��B�>� �.G�ѯ��2 OkَM\�3iM�;�Ƞ{�!�h��ү´5Hj�}�������I�F�,�&v��.�B�|�7XhL�@���Y^FUY�t����k��~`�[��/�j̊��ͤ��v����l���L�-���� 6����0ˋa]��ML�Kd��Փ�v��Y~�h�HV6�Hw��!0Fx����]�$���L�Ml	f���MQ����N��V�g5��Xn�h�R_�Ln��� w/*)��u�кT���ϕ�:n
�'*(���K��]Ĥ@��ǮK�������d����^��UZ~Ϣ3d����^(�guFmx,5����|b�{��Z�7@ވ��{�a�Y�J*�u�bpf1���R���"r����36��I�+�5��|Tr�=�,�0�L�Of�XA�����%�_�w4 �*�O��萤� ,-\B���Nnq8�W/�4�L��+U-q:��8�S�[װh}���[��X�6�}�a�:#��H��lV�&�2C� ��i���:y�l5��U9��Q�)�e�8=�h��Br2D���I��
Oӥ[6�zn�C��xf��E�Ҿ�����ǟ W2a0.�L��R�i��J���5����d�>8)v�#�4 �LJ��R�T���r�p��B��Ƒztm�"a]�(]�$�o��eݭ���?M���ޔh���qᡱ�'xY�S�$}��'.��H @	h��mx�%�ג��5�ۣbY�N��x�э�̵��N�<��֡~2 ��a��B��}�`ɂ�o�ю�} ����[�7�*���P	���o$tU�bN�*!S�KU���y�	,9蒁v���"�K�C��9�!DT�'���*��G)s�Ɔ6��8#������vW�l ��uV�`�sV��|���E@�%��&�@�}?�q�%�=�����o+}(%ӎ��� j��Y�o㹖;�[ ��(!	3r����>8k��Lߐȹ�*��T |�ŉ�.�����f��U �h��bC\�(�����	��P�+q�Gߎxn��j���i�33�T��]XP������5�
�v��&Þ7W���c`^|M6K����a��l֊�� �Y�0!ŉ@�Hu�:��5%FPn��l�VK��@lZ;S���g$"��!���'?�f�`'�Z�4�f�u;uC߅����41�R�.ҝ$4f�@e�ﻋ�dO����������{+���Q���Lm�Fr�E��Eݍ�+f����ߟ�6�껟�B.�V�Z*4o�馽��X�x�*>���\,p��m�����b4���.�0Y��������m O��B�!m�LE���#J��E�\�ڭ^�;�L���������p��W��Rv-�
������:�Sۙfz���Rv���8φTZ�ݝ؀����K���`*���WJ�W����^��Л���� ������	h�uQ8_'��ʩ<U��sլ�@Q��tQ��Ά�ӭ!�ݖ3�k��:ﶯL����f�`���ف�@�����9x�B�����ZuWa�RԶ���S�&���}�/�ʧ�r[�W��)Ԝ_=�_�� m@ֽs�R�ְ�ab�������z<�9U4�q�<�d��Q�m�l�z?�����4H��I������^����x���o�B
'M�&MX������G�˝v�y�&��FMkgƬ�ʧ��w?�u��M��k;�vHj�"��g�'�� ��Z����ej	��n�l�:�9H�A���%�7�3����;��-��

��V�m.Xj����1���ѣ,�'�Ӈ�	o����Xn�Q�=�_=����&���]&�8�2<8#����Vl4&Y���{aC��g�i�o��=p$���>���_E��r�D�}�����<����.%<Yi�w��{���.G\	?�_��KŠ�݅�e�@�q���7sp���<�p���F��0��s0.���4h+�]����-�X�D*;�y"ZZM�l�SB��?������;�1��c�C�t�`	Ǔ�%[�T�F95M�n_,�
�K������qħo+�Q�)��~8e(��+��`^�����������
?GliW�d�� �'��1�S:X^}��y�TF�]G6"d���K��rX���nǛ����~shv�Z�K% �]!x\�"ϔzt���҃��a�_j�(msK��>�Us��#l���� ,޹�H�e�o�T�5�����}����L�-�5����ҙ��W�)���A��Xc�u��"��V�(�K�D�T�Ҥ�ވ��$���C��x�w[#ݽ��+�q�!W��O@�^�| �� �]�Y��%3�¯�9�D��dGP,sk]�Xƫ�`E���1�cCvf�W ����"M)|��fVW��1�U���U��T�^Ue����>3���]����kH�T���XcN�xLP'�y�S��U���r�끠�Rt~��8Ym���Nv���\����U1(�����m�O�`��O��f�̿�����C��!'$@8�Q�_����[;OӺ��>j��p�ԃ��$��/-N@�]��W��jET�OK����?KtP��F�A��N�5����0���o�PW��9Z�����:H=�&-R���u� lg����e[�Y����u���n��5��n���}{�~'%��(p�Hm�U�Ix�F|�-R�!9���j����]*=� >7=M�M�~��q�<ͰW���zߴ��d?�+��@��f�����+G�v�g' F��G�ݞ��q��b)\��o5��{�u���N9D�}pޑ��M�%vE����v��"IN�'�������R�<�E5�Tj"�f�3}EdÝ@Cǘ���Eތ�E�!��%hsm�
�װ�yOW����`GWM���j�x�q�#��������kL˼� ����"��\��k�1����pY'XA���Cv�I��������çG�\�X�?Nv�%�/]���
����&�iy҅Wc�8��s��Ⓟ�ƻ�WN���`�x�Qҟ�S�T�{G�φĦ|�J1�E�#�)y�����~>��V$f�g�ϒ��o�0���>@?
&)c�sө�1μ�+��c){��/��1��r�Z?�l�WS��R6����blk����:^(�����M�;��YwQ|����Uׁ����3hO�_�)o�o���<�� �ʊ7�a@%i������w�B��)x<���F���](��(S&�)�bmS$`�x	DI�{/ׯ���ꮮ�$��I� PMӇ��@$?p7�<�]��.���Qz�9�`��x�)��Qm�L��kB��q�'�Y���\9�#v���y����҃��)V���)�6�?�c"����+�K�&!T���A.Y����3�W�Ӓ���J�����uu�o�h�_���]1)X-hJ��Z0�V}��|���� ໱��-��m���w��&��9���e�N�bRq3��ox�*H�_]����kW�[�Tq�U�|��B�&�>ٵu��W\cq���#} j:�:�]m���%���*�2Z�z�����IL�n�5KGZ/�EU>�[ȡi
	,hX��qr輋xZ�2�\���.��b^���-s�"��̽��v.W�?���?�zs��/)ð�$Av���b7QS�ǳ�<���b��?���Y�[��#������$q磡�?:��}���2zC��]����������Lu�\Q�R��~�q��3�����Rs�LNtClV1�>�I�ϰ��k+��:�431�6Q�8du��O���)+��R��|9]�RD��^�MaD�G���uw#q~�,��3�ҭ�bH���[Gu�����3���(m����LJ/8wf2V=�Ю9I��%���b7����1ڂ�����!��*�=l�_�n?��ؖ?���LuF�[x��>�bmZ�M$/M����}}|T��Oݭ�uL���:ppS:�*���in�8KN��';It�8�b�ݾ�i�;�E�1��<��z�l���