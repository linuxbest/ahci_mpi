XlxV64EB    1841     880m0#�:��x���	��ڲŤ�C�
A�|�b)QRЛ���P����SS��J"R$�%trgy.+��\Ur9�vU4&O��OSC�~�@c�ȳ��h"�T�f 颂�*�S΀�ַ;S�:Y.mā���?NR���L�RI�o��k�T�=z���W�LD�ֈLt�~Tp�UC��µ��R.�$�����`�@���!h�h�rV�����r���,��m����~r܋��C@#B�}�{ްU�9�����`�7��󬖃~���$��H���b!oI��x�ѡ]�#���H��H���� W�e��f�!ZQ&��M}�G��5��ү:Q����G�ۤAj���}jf���#��p�Ľ���	�zX�Hy��g
���K���5?9�2�A6�2𞸚
mF�B6y���W%�4Q&�����V���F�!�uo2�����x�Bm*Pt�I�D��G��Co��������ٟ�]mZ�P$^�g(�Ъ
�[d"�/�bL�T�Y����"��u��3ayj=�aG�>�a�e�T�q&4m���$����vw��ܓg�!eU��Ƭ|=u�qӇƵR�wX#�����ĝ��v7���L,ڮ�<eh�|�g"��ؚ��ˡ>�r��'W`�W� �����\��q�K������u$��˓�W����D�o���@K�� ��w�c�G�Q�G���&�Zw����Ƽ�S�ïE��W@\j'j5K������N��R�#�2&�V�����9Bs~.�PkZ���=Ԕ-�X�^�1x�l2"HmW��oK_�9������3?tc�r㡶��de�˞}�%������
�u��k{a�#��0 �D*Y?�B��M�#�)H��������&{���jR�|�.�e8='T�ɀ�UhH*���VH�[������Vw��A��U`�_���Ph��y��?u�%��~�<��6yО���O�R�~f<��ͤc�u�'��ԲU�d���K��q"�õprWl�X�P��ע�Ac�����*�S��'y5b�G�I[!톴9��ܽ����aJ��5>�|��ڦŧ9'��e�r��Q)�#X\�if@?0r@�ҵ��ѤXrأ�sV�T�Y
��\E�g32:�"�����J
�+����{AY-�2Ȏ�������#KS�s��lZoL��jj�<�%f�uݳ�?}���?�6������	3�W�E��}�Yi�?��dl����ڮ'�����f,��%��z�iG�-R�|%͉��{E�pp�~�N�}󖷏��(�(P:F�'-{i�XNNx��@����.D~�=!M�����w>���R����v�L����;�K�3��z���J�k���M[ծ��_v������j�l�Y�����e�B�|�5�n�n�:�+\W�xD�㠫FgD�`_ñ3k�U�eG@�8����Ӱ��ӫ�,9F�8�܂)Xh��u��� �W�P��[�CǮ�Uu0I��4ɀB����qE߼����$:���l`�Sw��틖�d�$�FV-l[Vc�!���YX�0�ȞP��vըD~��&�"H��tg��ؖͯ�������UK{w	��s�;�8�ۡrФR�$�Rx�����H�	�N�ĉ9�ϫ��ͭ�T���_ZA¥�/�`4ޏ	<��NY��E	9$��K�I-ߧ�x���v��6�ု}��g)�+�$ݑV<!�����0זW�o2P���ڲ��,Xag��RjZ����J���Z^�
%_�R�N4&��^ǈ��蠓��T�C'�mAKZ��8�zq���*�6E�~c��嚫8C(�1�{���8���Ɂ|�Pb)W�J�����E�B�	cMu�㇈x!W�鬆�<�H���˒�2�+SJ5�:��U��o���Ռxi#$�(���n�k.>U�9)i���ӵ��d�ϗO��I��P	&y_�Mn��4�7J`�w��*&�|J��8��ox�@��5X��17�qvZ�NH;������8����R5�,Q%� 7t����,f�g��_&�Hi��s9� P��:0_�s�!��l��B�)2�3G��O#�
IpvO�j���I�{�`����)�ur���M4��٘����-�[CLr�8d��~mz����j�.�8��U