XlxV64EB    2e1c     d30p�@�{�+Ng,\����#�yR�i.�.�D�L~R�ۋY�`�������Q���6l�zCK�	Z2;�n�3�	�}���"S.�e8��$c�N�8�ؽ^���3���fV��)�	�L@'@K9���s��$�P8�T�a�C9�z�N�S��)�t�W��)��:�^��k�&MC�4g�(�c���\Sڮ+��\��[0�;�2�NƪQ���/v_4t��ơ��Q�gq��{�~��3�a!�VY�W�myk�Ip��@���B̰Mܱ���}lr�������!ػt��S���ȗ>U*������5q�V�T�Ӝ�|W���.�2�Ti�u>�t��|�+Px��=oFL>C��(s+�H]���!��N�b�iY.m?ʲ����7���b[/��4iGIR�k0�ꆭ�,������ZY�B^1���O��<���'މ�Br��b�v�7������ҟQQ-�}~h"� =wC2���z� w��vP=���[�W�=$b`���@���`ӦO�1�g�O+�g�ړ�=x_�h$��Z/��L��� ��L��BS��g�U�Z�~5Y��+;�&�'��Vϝd`\��!�Xe���-4�˘��o*s�ԋkb�"9�_x��ב�T�UnH)���k�N˭�M���g���|�u��<8=>��ц��̋�
�E�I��$��>r�Z�$�cFp��d�̺�E���](.�B* ���1�}b�0�F�nف��֦�ˊ+�h�'��������Hr����輦�*�OLD�>A����N�1�%Jr��U��nHND͢��s5�� ����1�rˉ�
_�w�{��{򂾿�t�*�049RI�e��}������y����/n��_���*1rƕ������lm�ȣ��y �J�0�M� �5^�wݚ�t��.��GG�b4�(�1�=i��	?��_�I�fUd�fi����_V��{���`+�[��?�bO��wD�2~�:��qZ�f��a!=!P�(�v��Pq��Ϭ-m�=��Q1P�Q~�|�ç�c)e�l��������3��kØ0ˬ<�d&���w�@S��?kC]��L__�g�kDWc� 4�A�@�p�t����4�{�0���Wz}$m+�>j��h&�)��%��F�X�T`�r�T%�B��G����Z��Sd�Y�Ö:ɚn�ʞ<^%�X�~p?#������f�tY���Lm���s�5P�x(�e���y1�*	s'^�G�v���d8��K!���;����db��i��r�����Gږ��p�������٥�'qQ��c��甮�p�|��y�6�0�U�
�7A9��, �JL�A?X+ڡo���s9�J0~���,8�����jy[
P�Ϝ�,��q�EO*eP�l�5���G�$��&O�89π,�gĊ����D]�ә@��E!v���mצ��+��\f�ގf����$� �旴�J�͈�������A�!�=Cq����L����>'U	�j�@��-���Vw�`�w[��/-:A5٭�cC~��y��y8��D��p-	�m
lZ��-j\-�� 
�Sd�4���'$��B���]4�g�+^�1��&Y���H�����Ⴇ��]��M>v]6�m�m&�%�ܙ������O�Z���J�pK�2�T���!;Nܫ>5W>�e�Ϳ	�.|��
p�z��_Y�D��SIfR���cC�'Ú�f:�]��n�IMi���R[[�P�\!'��)�z�����Ԥ�/a��|P��O�Ru�Պ*��6N2�)�p��_��ŽFGTA��*˶�x*!��w�EN�:^�M�QX����t�5Wz��!�*�m��}����TU���	�sܒR�� ��v�gNǲ�xhM�\!�\njD/V ��i�����xc��`��/�y->�{���YP7q`p%�jy3r+�Z�����m��w��J	u�&ZX���=��#�B-S�lX�x-�U�Tv��|�7xING�݂.j����.87/���S�+�G����z�KY�c?ͺv���������K)�!y<�t	��j�ŀ�k��j���r$�r ]��J�r4a)����W���U)?h���O����l��$/�����s[�*D�մ�c�m1B�Ec���(��}j\�$0��*gY`�~���:�ź)W�C,G>�/QΖ	w!����3֟laj4�&�R��+��C�9�֫堕�K&@h���M��Z��[�j6�3�Iy�C�$ Z�:�3pk��$��U��+��- ���\'�T�Bl��g�$�]�����Sƅ�����}Gh�5%�0����cO�B����p��&��G3=����U��D�Z�!���Nh�3���ʣ�sT�vAw��[&��l=b�UPh�Tя+�OB�6�Gn�Є�_�?ҫ*D�ҹ�SC 
��B�uawەQ�H2�����>S�|���d���f:�(w��I>��;Qֿ�`��eS�1�¨�SK�~�%Yx:hn����`x�oy��F�� EzZ��B8�e5���6u��\y*����Q��*���i׾j�ۯ��uvX7���R��#�Z��3��6�<�Y�I�c~�lR���vO]�'��˒6�2A>~G,Q>����ģ䀭)�:�;V�=��or�������hh���
;;d�BD#rp���XB(D��a�]]q���fÙ�NSQW��:�g[�w���R
t'�Z��2��Tq6�Iµ��"��W^ڤXd*s��W�C�����3��O����S��l��]�TXt���Xc�~�?vx)|f����4ջ�U��-ڣyt��֋^O��Z�A�j��$��N��q��R]��\!u�Q��f�Ĭ�h��>g��W��F�B�y�࣊E#�i�y=�)P�T�=`�V�~�λ :.����Ǫ��7s\�vMƲ�L��՞I�3�O�r��#�K�|E"dw]L�G��<�Gݎ���!jc������̙�d�-�J���KZ���}J��W֜q�����/
�17^b����M�>�J���@�f��Q�&�'��cLB�n�������H���A�[��-rqBG�eC[5����׺�of}�F:B�ǣ_
�1#�z}<��N�i�	Y�/Xu�b�96�	��ʋ(e�NX�^S�QX�	��|Ҥ�_({5�8����%��FT&+H�ʱ�f {j`�N���ky~�t������Dsd�\t�j5�KMV�p23��߂�kY���`�<R��e7���>�<&"�Qɩl�%����0���|�|�x����:����K��[����A�h