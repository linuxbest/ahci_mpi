XlxV64EB    8a3c    1890�~���)�k�<�����?8�Bf���*�����E�R����#�t���4�I��A
�p5�)���R�'o?\��Y��H��Gk�9�.�ט��qI��*{k���j�z��j��
G$^w��&)�? �◰>��&��8m�-T��u���n{Nc&%b.�)��\*yb�8�7�V ����e��� 9Na!���#x���܉%{C"|��U���9ݥu�tl<Sna�@e���oX"�w5h�e'�pC��$Z��;$l�:kD纨���}3ҟ��&b�!֔�ũ��]�s�Cl��sV�B�R9���8���:�ۃ���i�:<�S��N�:�ה��&����<��M0�w��Ƚ�Tʋ�|&� ��1v
���O��٣LnkT�j��#�~2�%]�o��\�&?�e�2��*Վ`*��h���F�ZJ� �]���E�ˀu�(\���udV��-CDk��XåX���!�hi_p�9�.�Jv6���K��h�s��3�2b"~C�0�I
3�A��I�W�a[l�l���+���ֱ��<ĕ`�δ�@��ȚѼ�z�8�ʐ��&��┛��H)A)ߟeԻX�xV:�ڵީ]��������u+#�'	�dg�=\@���T����?m�~�&D�į��\Q�C��Fa�2(�u�'������Q[/9�GM���D��)G��͠���$B��R%nV�P� �6Fm������G��RM�j�"x�x4�W�w��F�<����%��q2�ȨߕC��	�ǵf�$��}h���ؿ�G`"MZ�J��p��ݶ�a� `�	}~�aA����K���VY�<9����P[�9��` O!�-��ej`.)�CE�{�#V�$�Q�!zr/_d�91b֝�R���A�g�e�]�=:	�&�4ǝm���c=D��j��f�y�r������fu�� (V� m���d,��Q�Vk}�8���C6�d�8:fg'�*�eV�LtxiC+W��]'@�?�v�`�A�ÜW����4�\���]�.̫�?��w�G���S�u(�ί�͑Ȫ�}F'�����;�ZKڶC�9�i�J��٪Z�G��YĎ>`�av���)&�ѥ����g�PY����K�b�����)�c��`}��gA���Ols�+��娟��U�E8p&�h�ݒA�jͽ��0�--��lb_��n���
�R3���FӰ$�y��%��`���&'��j���m.\|��l��ld������B]�8yY�^��?2��UM��J�a�Q����b3j�v�p���/��2L�2����v���RO�pn���D� p=������_���A�팫E��@��:�K'�2�'Dn,^����sHMD�/<�)�Uej0�«xMU��0aI���>�DM������K�Qű2d��n�g%�y��K9V�M0Μz5�;c��s,k��̣��F�J���f�������$���38����k�}�;ͅ�[K��O�'<�<��]�}���������G����4G�����l����6ˌ�}+�j[�b�]�t�ڬT�h�����͂qF��g��	,t������{d���W����r�'�R{..�\�n1^��_{�~��P�pL�����q�]
�1by�
�(�7��*�~ש�� ]�<6:��;���Y��)��
\��1�(��(��[J8��Wg�⃈��eq)���S/���
~��?g��'��ط�(�źc��{|�%��ߠUP��0�㉈\f�^�F��8cH�ULAϥv3_�ڄ�������!8��hx�2�P�/�$')Ё�:|jr�4N~X�kLb	&EJ �_�]TU{Ho1/P AL�%�'*3�A�N��T]�ؽ��-Y��3'4ccmYH��#�쌿��pb��b��CN	�B9��?5�����8 -!�k�>���?���d��=c�}�����H��O����K)n��{�i�h���ϵ�>�j�è�l�*D����.��>S���珫��EE��1�hգ�]׶a�/:lH��Z1.�]�s͉�af� �
:R�D�\fYRwDaNq�� BFhUd���ط�p�S���X���8����o�TIEΈ�5�����9�i$��P�c�1ɂ��Y
�Jl0����3�`"��}��?OwT�C�Y,��]�ُ��kq' ��s���ͺ%�$3��S�͠ߕ"�l�&wF��X���6M�m��в�J�1����T�Ad���#���s����ݱx�Z3@��Kړ�U����~����J��3f�jim�.CX.�ax�_Fsx�6�[wL��anAp	�����0��}c�,�⦁�ο`~�̕g ��+�SN��?�4�ޘ���.�%�^�F�i1,H��dL��q�w��E���E�X��<L��*yƘ��p�z��,��rS\�Î��I
V�Y�DUc3�3uJ�jYPLc����>���pr�\��x/��Wi�m�9p[ By���{u��+�P��l�z��]���3��5�1"OIK�P	]n��kz�~���&����'��p��g��[b��iY̍�Բx�p��?��\"ʛ���/�ū#`�GI�����of͹ݡ�j|�b+�i@�������6�����$�	�Yr�`ţt��Ԣx?���>����ZD�^�f%*�g���D=v~��ǿ��s(^sw�ӥ�����k���Vǿh��[x;�<;tm��/Wu����ʯ����pa�"x��-�
�˵Q�f*����5_T[B��&�6�&���*z��ϐ#x��Z�����M �2�MG�&<�����A����2M��#�Y���V�*�8W��
p����_�����='�E�e�d��p�+�#��K,������H�<����I��4<��y�B�ӊ]�M����3����N��.a\�,�1-��"O�_��y�ޯb��7��^x�p�p�P�*���@2�I�a��&n����+B��>�m�c�������2���g��nJ��"xҰ������:��|C
�ˊ�5�y���P�����`��n�p��������h�>������0��{����bP��̮��zNUu�ҁ||rZu)`���\C�2�0��2���N��A����0r���:�b�G
L~�,0�!=#� �}�DN�P��A|�~Q������d�/��Ql� ^ӳ;�7�U���+F��*6ޅ�Hƣ�(#��������Kj��I�)�9�)=��@�����k�'�4�Z�����]
����o�Rѝ���A��C�(���Lc�0x9�Q���Q���Vx�J�
�pہ�fN�ʎ"P���?��|e�r�	/?�9�ޝ#����@t��������J��n�|���/�����j"u�
����.O��1�q�b�-G�g*�t(��*0��,Ϳ��{��{�&YcC�������]�-��U��U[)���_w�OQ����k�� �@�����9��=a7�H��Ε�w���"<���a*�TI��%]oO�N��J}�Ԋn���CKS��n��g�F�~!�5�{Egh]�7�6ld�L���;z����p�8��"4o8�7�T�w�m�4P�u��YH0�y�>�,<x 1�,��w#��gad=�Ů��� L�J��,�=�Vu�])6�ha�n��=��2�u�q�(�*;'{&������ݝ�O8���;� ��ȴ	�Vد�ؔ�@�Hh$0�/kbR�D�?-*�qZA&�}5"�AV��Э"##����t1WXS��gZi;��IlA_d�,~>��5�5|��!�h�8W�.;�	���7�g�E�h�1��ZԂ{�#�g�}옜.��)��[�ۖ�y&|Z͂$��#��2Rpg��;�\}&��	��jf�E��]a�r�p����o��3o���	�E���J��Ju[��jt1@��U�0�Gĸg���_^��GmҎTN�1 ����,n+��Wʮ���J���_@�}����p�� ���`:�LE�Ŷߋ�&�,��CE�-x�7�݂qQ��c�����Z{
�y���B	�Is�[��9g�2G��j0kB� 8V�{���+���=���Ў�ߟ>�m/�Y��`����V�:��;ɡ2v�-��g�q|q�B��Qm(h'��'7E���eRM�(�IY�^� b� �Җ]-���ԑ�,9�D�L&���|h=�zZ��>����\3�P�����1�ޣ
ƚ<pOl��=�u����R��f�t�E/m�3{m��b �����
J�`F ����?��5u�߫%|\�w�d$�I�^P¡~m!@t����?��0,����N� '�G�$d�}#T���.���t_��7;P3�|��@���8���K϶i�, �f��;���+�ٖG�+�q-����F���
�����ܖ���t�q�ۘ����M*zW�텵 ���]�%��|�%ܭGv�����s��W��z�����l6�g�ƚ�R����u�Ow��$Խ���!���yɟ�I(�R#WӐ�,J�XR��c)'�ҝT�+�z���ơ��8�Mx%8 ��ҧ�����G�+��zϑE�L_ݧ���fX�vĨ��ӂ�k��~S7iK��n�s�0�P�Y@N��3���|��x>7�uL�>��]�mW�&sk��Ry����ه]�P VR��Ybo8������N�Q/F�y>k��^����^�T3ϟRC�|N9.���&������t����!p�����P�r)wd�2�񤉦n��5ͪ逅�ph��� ���"��r��5���0�[�ͼ�㾋Y��^3"��Z��P��ەm�,�چ4�}�U%I��B���z��艠�V^�m��r��ޝ�X�9�����c� ~���:��W�x�4�Ҥw^��M�LM���\J�������A��^`Z��6'B'\����Ǆ�,o��4�5� ��Ó��#�  M�X���-W��Lv������h7:hE��� ��g$����ה�
�\�ɑ�w�d��x�qG�75�Р
WUҼ�Rʱ����߱��k$���>�o�9��V*3��V�WV���LV����2�fx�*}���RU0{h�F��'�.�淚��C�?;��՝LrD������x3�Q�6@x���k��둠�˧�����XP5E���1�pE<0��/]T3�8,@�:Ć{IP2�ǧb�Q}�s˯��-�Z�>�p�r��{$3s���f���� 0g~�|;&,�H�& ��Mޗ�p~L��AE�6�y�~b��`��yI�g�{x7wD�Wr��s���X`��+������5w��ac~ޘ�>M(���=�y���6��6�;�󮵋��"�I��:�-��hB֠�f�ͺ��yIJ�+�7�^��y�:"��ù�ޑ5�˦���=�d���>wY�8W٠\h)����^�2�10��F;�I&�Q�X�����ho��1jig�.k�G��1��4��s��J]�M�
�_�J�UՠQ`�!��f��<�a֕�N#+$��D�������MGNg��%��*U|:b2�{�D��RT�Z?�a�N��5!���o~>�=��H"�ZVu�w��"L ���l-�����k�����~>��i��lˡ^��]8k~�Ե�*;o9���P���6�'NT�L(7�~�gNL��1=ϢD6��H�i쿗 k���[n?�ܮ>R�&vlG��`��j��?��qɛ�e��4�U0 �ϰ�#�]0?���Jf��a�z����`�1KXy�d1g£�p��Y��4"�㘘Ͷ(c;�K�7����k��Ս�A���p>V��+�@��v��&΄a't�������R�M�t������͔�D��%��|kM8S`2 �* �Ђh�#�W�y3�5��r˖(�\���[H��s���g���Ĵ�6�����i����� ��F	!�nxd
~?�Pu��g�h�U!td�ޥ�s��6>_p�6Q|�����׉�'�#����T\r�	��u��VwD0���v8�<��hs���交"hVqn��d.d�Ǧ`Â��������Z�5H�z�#/Γ���U��ܵ֪��t�)�;��4�{�)�Q���Q҂�%�fX$c�-��m��)�����+���L�aP�mx