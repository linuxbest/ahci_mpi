XlxV64EB    7100    1720-��D����٭���#���VF�%�gi�P|�ΤV�D6�ŏ"Cj���������U�˶�5����ٮcB���~a͙˝Oc�p�<D�M�Ɔ��B�K�^&�S	�dd7ts&�A�F}YN0qu�sa$�ި^j}SQ��+�I���s|����`��$�Qj�\��lI�H	�����"�QB7��D�è1Iû�w[��.��E0��O�҃�f"�K�(�Z�#L��u�L�$�
�_$��5���E�hT��.o����4�T[v�i���������R��D�Zu��M�p� 3z�Nu^��xtO���O#��G��;���U�Qx���!$��C'7�����XWGO��NM����a�d�H�g��d�CZ�6% t�x�O���z��u��C�	���`�"W�RQ��I���T����W�v�wU�ld������H�,�{KD/�*��YȗD��[̷@0�^�Z �6H����c�,x*����% vg���mJՇ�"zb���=�+$�Е���ݞ��3�"���{P�M�<��3w�_F�P�KRǆ�A�����4Lc�lt����2�s�S.���EϨ�*�\혟��`��J�����r$�E"[��̼���%�HsUͿ�n>M#k��}�j��G��;$��)�b#N��ܻ�����{�D	-���~6�{�k��{�@�R�؇K�!R��T���a���!�Ʀ1�RLVn�č �;)���A�w���䀰��s/��;��4�7yS�o�����H󜽙/�{\,�λZw�?"^�6R���-{�%SI��d�&W��O\$��K�Vx�
��sn��2�NG��疁���e�DN��Ŋ�8}fOm$�����Fȯ�.����Z�t�'�`<Mt���hE���02���qm��AR�l�����8FES�����؋(_'v�;�����M����p�Pa�o�z����Z����4��|�����|�*2��}J��r*o���V�R{�4s�~�*k�ډ��� /s�!��ہ��*�N�es�����ܷ�Y� H�[���N;�n{N@��/��)'/$H��#̃;"�-��o����������#��:�'�h�Ad�`{$���G��2ٽ�+�b��&~<Ḷ$�ta:+�pqI�';�.���Gc�*|V|(B�����[~n���w��'��
?�;֨g���<|�D��+�-xp�U0��?�si7�2.(��� -���=!d6$In��~X�2�V;�LV���N@ӹ.^<~e�eG�z�Væ~�d�'�!�3��*��C�t�Y��BTQ��,Ǐ�)����sR}`<b���P�pD�\��ȭ�Y�*pw�[2;����;�. �0��dg�R�l��&�u�X�dP��\�����ż��ѱ��S%u���8>Bų�{����D�l�̐��%��$�<K�Z]&��(��yҍH��F�F��
�b���m����yP;�M{;p�, ؟��m\�
+��c�"�T�
�o�t��M�H���bY�'����pR�OZ�S*JL`款�f�[ˤ��R����c>�-t��S��Љr��(�cR
����A�`s�����~C���c�cv�s'e�M�+%��8��A!������	���$����<�Г�Z�mp?R
	ׄ��_PfQ�z����=�Pz,�u"(Ũ?a�2�Jm �ii��:~@���>��D�X�P�Y�F�"�)���A�z8h4P1F}T�[�qo�� .l��>��c"�i{�X71�A����kŏ��4��P/�dfc'7˵�C���=`$L�h�����k�Y@��胲��f�gnA���pUI�ϲ�Hm�� ڽ5�,�p�����yj���H��Y?��.���e
{��s�:�(*��*3R��C�Zp�n7_���c>�G��ө�=D.�V%�?C=�/W�Kz���fr�=�E����`doa��]�	q�?��s�!�M��,��W��@9��U��q}�j ?�Ly�劣��՝7*@Y]+�+[�١�![�\�D4,�B�́���j ��0�w�g����X�v.Y������z<��Hѥ�?���v0���)���0� Z���}������*!>��z�eǐ4�-ŚS����a����P��sUv�C�U���nBdDe���g~��)-1�&K��6��"��6�Ⱥ�sB������W�m&'�K�טx+�?#�����x���M#}�Vf���Y��o���D�#m�/_'��/ac0b�{��"�qB�D�ˣ-y)�l[�xH"��ㄛ�)���2�jAFl��Q0�����y̪"�w�.B,5�Ԯ��o|+��s&zn"��B5"'�2uб_+���}4{�K���Ⱥ3���Rٙ�@t^��[녘$��ùM��cqf�3}�;R��8�ݪ=�8�=c~ Uz���a���:���rU��-Ґp�]|d�><���"�n]�+�xN��&4�O=���c3��/�����T��Qm*�Iq��m��w�$�8��>dNE:YA����m��2��h}����30�@�Pq��� �z�}&i�*Zvci�����$���e�'�6	�k`�J��]8��1M��C`����H�~�Js��0��Y����g��ca��ցY�X����t����E���ݟSZ��H`�wESA�&˟Lk���5���ː�L��̀���\"}2�WE�:�q	|PM~fx�e�nPN�:�tS>��Ƀy��� �C�,�G�On%������Ϸs`�C>v��W����!��q1J����Q��0��	mSe�:x����?��Ls7��K�2"�K�7m��� v���iU�-��&�f�ƣ�Ծ�Ko�3�$�i;]D)�k�h�b���"����4����_���PR��_G�ԠA�ʎ�X��`y�Va[�����gK(�g�jg��VB���XT����Z�����t<�3�꼻P��7wI���~+�"�涧.�k}��Ug�@�.�Dٱ�����:NƗ2�
��ʜ�JK'������y��<�~&U��뭩<���1R�j�y/GM8ߎ�ok�hX��� ��"��/�x��9K���会+�#�0���S3�_R&����N�	8�Η-c2�|����*Lr��ikn!�4�ӼcОh�������p�?23�`����!�x��`v�8|P糁��V�)ZD��,�8_�&�^��m�hc��e:�jl(k��|��k}ψ�~�|7kӀ�P�����f4X뜑�h�Z�/-���M"��`q�[�;񢀋�߽Sw��M�*��D�\��8�/��P�ǼUL�(ݿj��]�G�Y��� 3IY��(���9a�c��ft�q�u�M���)�RCfz�IHjE}�C7���߸I���]%�~7D!#0��		q��d���T{��G�:U�N� ��)p���n�x�HdF�z_��
����;���R�Yb���nӽ���~$I���) ���;'��&��5	��%�ߵ	Ip���X#�<H6ř���#�.w��%��[pZ�3{��a�.|�<�r�W���1�#��%�/l �w�u�W��YU���q��~���މ�7 r��jF�	ݛH��(d�ξ�hC����IX9�+ݶnz��N�n	-�PA���%IE�N(�P��4�y�h*$����hތ���rRq�T�B��y����C��ƽ��:z��/bv_���.�̿{����*��R�Lr�P2��E�<�ߒ��:&����H�I�ݞ�4_@~k)s����,fBqAɘ`*qk�>�f�A�ɶ��h���-B��D?�p#4���S2w�#�*�B��C�yg���C\=�$�R�#b���S�:�[�n�H�C�)�y|�V�``�aFύ:m,���@��o�X�1�7E2ٱ	Hir+0�~Q1��\�2��u�i�Fм�v��eA3�t���W���K���ǀ��	�H'إ�~|_A��Y٘�U����Jص�����&e��6O��s�4sHO��S�m+�@�G5c6t��3����d�z���&ѓ�R���V%�8��f�����f�S�c�(� es=9Z'�K:f�6}ZE��79w�"���	�5/�}������Ǵ���z�����$b�̟g��S���<U[Y��ust�*��7_j����A�>�	W�ɣE�O,��#��6�Wt)�ϵ����E?0�Cy�չ�����s��"��VI��}����7��w|��4%LZ�)y�/J��#�r52f�m��ɩxF���qY%�xm�-�:���3C�n]X�@���j���)��~��a��C)�f�h���|i�i-sV�	��.���@ү�vްyM6�[���p
���H�g��N�K�+>|�L�2Z�mi�C�;��A#�_5-���c���h����=Ks`+���i譅nYoh �%�����h�a<bՎ�v#�+���:;
��p�h�d�';�.XG�S����RZˇ�����Ѹ?K�5�@%קY����,�΄����_�@��l���e(w�5l� �w�x0���=�1?2�,H�SrE�o�@bvTaF��(*0����}n}(�m«SJ��v�%����2L%��O����������#}V�b�9�������@�?N�Z��DOW����	�s�w��߶��dԉ��.��<���M��.f	�X[%L�N�w���H�h�`��c���i�xT�E�VG�4�'��'x�73xզ"�Qa�W���`�p&M���tO���n�q���!�b�

��jS"p�v�z�O,�H���|݅X���mbNڈ�������������5O$���ĝC(��2g3>n!�Mی��	, �N��Q��5L<��Q�E��o"�t����$�w��~F���%o�(⤥ؗ|��5vs�L挝Z�Y�r@��
_��S9/w��%;h�]�����bڤ(�_`9�j�π�P���l;��[p.[J�piy�=��Ou{��)���4ܥn�6�Ŵ��&�����Q���g����W��9 *����)�����־Ne����۔����[I�4z N�X4-���Fһ �ۼ�3s�CrM�9�L�X˜�m#Z=���u'�R!���hG'�&La��.1��=7��5
%@ì2.}2m��@B0���{�̱&�|=�H��|������*+���뎇�`�F��T�q��㱎�xB�=|3�%t��Z�Z�5,Q�$埘���Ov�`K{��(Mv����%j������O�FS��:*�|������]#6�in��>v���w�¬	�$�62�t���[-#,C��p����ٽFv�O�!m���)�U��IX�(��v.7p����`��Z��F�U�t��bxɇQo�C�|�ƹ-MzM��Ǯ��}���£�$��qY���(��>�݈�G�ӹ���58�t7�?��,ƈhr懂0Y{�|��Z�e���c(�f��������+�%q�j?�t:�<����9�jq�ʢʹ���]JzE���� \��=�)~�=�-��[���k����Tx��������H��[sO��6�����g2��{�u��2|��Qhy��J��Ϥ���,�Íſ�r�oñ�X^f���&b�W	O��Hd�3�)s������<fSo`hK���f�	%�\��h�c`!7?k�,
PA��G����b|:_��}A��ԬݾVN�R��z�J� ����Z�,~���\�I<~���y=R�M�]����3Z[\�`��`_��J_������