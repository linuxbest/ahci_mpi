XlxV64EB    c9f4    1a50�a�V�	ד;u�� h�]0�+�AB�43G5o��fx��#�02 Q�{����8��
t-�����6Di!�P ���S�9�*�S��i�!��Z�Tf]��U+ZaY�_)�j����J��G��z+WQ����ŗ[��}nt%0d�!U�!x���D����r�Y�Ť{"P����L����l
���e�����p�_�hCV.Ը�+��T�4��FnJ����P8 ȌW����]�rr��b�ԟ>�R%��x&��BtO6P�d��>�����
������n��;� �H��CA�uYL�+d$Q�ݼI����NUj�=�80�J+R)�ܩU��3�(��N�i v@�ŝ,[��Ë-:ۀ�V��y�Ʃ�v��o�Oj�7S��?;��7�m�{�޳Z��;U�"�K3���Kݑڡ,�܎��i/���1ED
�_���s� �a_��c-���[�e\�2	B�&������8bUKF��>(X�@�!���z��,��(�d��Q,�cEnJ*�
�r�K-1R�qr�	�( �z��(�'iyCq��l{���ά����\f�3�+��^\�)�z�>i�k*�H�ܸ'P٧�(�uР��Xd��@Sf����<� >�������~�p��9���Sg�k�����bR3�����+��� ��ڪ:)����=5�u��=ΦL|!B�`A�Ua�T*X%�ĉ��[o̽?,XC�!:Ԩ-�|�u���<�Yoʈ?|���R+G����P��H������2t��$e�]����;�}5{�딩��S	��JP�X�3����<ڮ�"�q�fr�:5�������ʧ~ӆ �U,� (�h��n�:��_�u]�OQ�1�����$��ҷR)EkSE��]F�ܗ���'t��A�����r
��$�O���۟�뤙�M�ձjdC- +U��Yڍc5\�����0�+OƳ\k-�5zDQ�P�{�����=�R�ᶙ�do7K�%4�b�W�A�P��W2��=���?�w?�6L?;���I�r��&e�I��d�@� �����E}�h�k2�b����z�4���Z���ޜ��>U�΢Z����	d.���;�Y�̠�dx���m�Y�����r�^<@a�g!�z����X�|����y�u� ��P�8v�ْ�	?p���6�M
�����g�.���=y��x���l�C�|C�	{����H;#�8w�p�w��X4���D-ղv!qɋ��P���3�B#������S.�|� �3w�a�zzy��TW��o��iK�S0mY��Xc{S�[��M{b�t3:���^��vD� �.++�~�D��(�ɗ�I:f^!���kv�� �#��,������
���@��a7����hڶ�~yɳ����,�S^���	'b̕�D�k�x�q�@�4k�~��z�`�§��=��5����)���s�h����FT)����A�`���h����~cT�}֊]�(|u��z��I���gN��zaSS������]|���^��U�k+:S�HX։�1���D[��=�J󒢇����G]��Nw��wv(<	��a���Ozmѵr<+{�Iǁ
����	�=�τM�o�;Ī h���@w�<���wOm�7ަ� �>�<��D��n�p$�i����l�A�=�+�zF[�'��&���~K��2�~���� �]T�Vh>+6���E#�A2 $ת}� rFaeFg���p���j���ǭ�kwǻ@u���E������8}eR߶_���cQ��k+
/��u��o'c����������q�P;<��D�"��3
��;<�=�*?��u滣5���{T�Ч��z���|@1�(��~��� ���m{��p$Z���p��#�����L^b��؇���/Vy��@{�n<����-�8�K!'�#}Ŧ��U`��$�G+&mx�[Q+��/ ���",�tt�P����)��5���_�y��m(�DN�β��;��YK�T����#a����0�����qu�χ�3���+L"���]��	�0~�@��D��ϰ�����:��߅��\�Th���.�����{XHW��qP�I!�m���@Ep��<x05�#�o�EK��"骑�����V�^{�hX�خ'l�j�;í�S�xw��K:�ƊtK��_R���we�ۧ�(o�L#i�
}}�3:SH����[Z8���=�	�qF�n} ���<,ur�U�O��=��K�ԥp��j��\c���!P原1��K��d�A*��tY�=��:��6u4˵��im���b�Yz���B��_h1���wjZ � �$��{YC>6��J�u�)��{�xv.�S��Ȝ�5	
߄a��A]�ۏ���J������7`�	_t^K��;j��R���ΩN������\�kN���}�%�%��Ⱦ�0�J�n�ӞF��
�F���}&$��slE���8�������j	Ұ�#���9��
R�E;a,e_[��Y�Hpu׾4�\��f��!���<ٚ��T�֥�po�;�l�l�S0��3'�5��K8&�wu��P#=(�N���1���,����׵$��Y����^zO:�|�Ł�.X�΄0��j��X�¶��S*2H�(-q�(�2v�� ꥁUab��tf6���l�{�X�����KMV��$�c�����"�ǓcK����8���ktBd+�����"�ID��N�7�V!\��弦���m
W��L���GG�|d݈�2ӽC��:�2�����¨Ȩb0d��𤞯�'���	���e53`}x�
����'�[��gF�Aȼ�'7a�������
���>V=c؅�&lok�.C|+Ss�A�`YsL�G��bg!1�!HM��xv�V�8a�|˼ӷ��A��㨟@rø�{k����z)���9�3 >E�_�pC(N��θW���k>:j���h3K4ĳ�D�&b����#M�p�p�\�o�Ԡav��D8�άN����Dt��Ic%�VztbFͮq�u S��V,���9�HC��_��Ej������Xm��Z��!�9��_�5�Nˑ�I�{��BG�%��5�u��������q�Ȏ�q����
#M�2�Y��Kf�e�卮8��'��#��k!F� �e0�,Z�e����[4 ޫ$d��޹�t�xV]�z
����&�m����L˒��1�s[T�ԏ���f{ќq�A^qtNSbN����[KV��L`P������^.ۻ���a��^-�92��5�O$�6������u��w(�Ⱉ'��J��]���brpu�,��*4AM4��щ��}6!�p�+�tZ�Hnߦ/�_�!�¨�i�>��D�V�a�`%�V�;�u��Г���:��&�$�l:��@u�#Ϝd�N���$��
���V���0z/p9��C�a��ÿD�d�rn��X���0�@�m�?�d����PM���.��W�kuH�
�$i��J��2��I)Ʉ�o@������"f�1�8Ks������Z����Y7[s�7�4����m�]��:����r�p�s�q���=��i��67wD�ٝ�\��_�S�\J�Bױ��s'�3m�@1�jcZ�f.�g���]CV)����f�~�t0��=3
h�"W��۪���A\�/ʮj@a��|�h^.i#�'�#� �t�u���͞�P�H�u����%��z�pk��l���擿�'ط�bF�06���5!?4�K�H��8�W*�1���|���A�O����¿J�FD�sh!��������\dpểࣜ}6�cL�� Jg��Ӑ.�򎈸��Ns�vD�Z���ĸٱ�O�C�:N��<z��#~j	6hq��,@����̃!� d�M���(�,�P;��kS��+o�[&W���
���� �kv�!Jͽ5>�o�VBNYؖ ���+��+�uk$dm0������j�N��04�*Sfw:_3N!�
��B���&i*��hm�I\����sS'Y�	J&�T��ȔH��\�����6P�Pm�g��u�|��[��K�4o������Id)١��g>`h��)��<W�ǳk�1eҴ4���Cc]���oN��ح��:$:"�A8AӣE1^Ⱥ�7h7?�k�E�iW׏�Pfs	6��3���E�1�US� `��K/��K[���F�3҃��B[�T�3M(�����8���2Cd�Ę-ǜE�k�Ķ��l�#բ�_��UV�f,�(�$	��M���S��у�gq��B ���<�y��VY�T���*aW����x|0��2�o�
}��P�sK�w�(�u/a�Kag��6՟���:3�k�P��w��.��c�i+\�cޫ�$�����IW9̗��~O�&7���w�1��F9�9�k�~��!m��������	�4 _)���ÿήDrM�T�)�H����E`Xʈ?��='��9#` l�x�r��Q^��S��Tي����KN��n�����T� ��E�@��L��W��0ס���������[c�����(�<C�-5��Xӏ�3+�����T�{��`�aV�NW��K ����/�������Ϟ��X�����z�J]�����S;�P����1%��`�H%-��N�&iݩ#����Du�!�Z���|�_=,�*�_}JHw�y?]�&�j�Ը�7(>����g��
沕�4<��ٍ{���!*�$��cB-c��:u�����0��d�ֻSD޺-R�'Y�Fm�<z�°��b���Ņݻ��!�%�#QU}��k/���4��;AR�=��F�f��S���ֺ6��ˋˑv����HR�YϩM��%�ݲ! �5Ŗ���L2J����Om��
���t���������픡��s��TB��B�*8,�����T8�s�΃���43�<�t�q-$�-��^]�>5��~6��)�)6���ɿ~�)��̑����Ϊ�܎�#�5�ϓk��TO��G:=��~�j|�����2ڒb��X)�o�����J*�9��R�	11�e0㯑	�L��ۑ�[�_Sa\�~��f��=�T2��;.)��9�8�ѱ��|=ma�X�JA�$E�ơ��4�`b�u3 )U��nA�C-�(��l�6`I����FP�p���&���?��y-�����~z�Fp��Q' b;�'�(�G�e�7m1�X����'_��Tu�B�e��ؖ(�}�������`�!��RD2��(h�cf��*Z��g�SF�3�w��A)�Z^�b��)�.�ƌ��0�3Q]/B�!�=��.j����# ]&�6����Zw����Kg��KL�Qg��E%0��P�/��&c��u�gg���7�͸K�HEc���mxj0���8+�`�E�=î��W>m]��`����}E@�
���*����re'����d�cIyfKOE%�x�Á_�ud�)�2յ����9��bJ>	����C�`���-��8�h �=J�{i5U8cevz8�2����$�i���L��}��`�����$���d;V~�f"sUrf�l����)�{_�� ������W5��tߗ��̤��s�IGO%Y��Sk��a�O�M���e�����9�,���,*�@֊�0�I]giYr�p)��%��r��V�^t�7��/�f*tl�;
%_ j!6SɢE֯�ϔ��5�չ��[�9�����\p��g&�9F�xbP�	�����S���3��>������_�C�����g�I�\{n����@n4x����Om�։�9�*��J<,���k���t�D���tKb^���yv�oג����E�P3�n����n�}�'[�#zW�I���e���&��i.�s_�����Gv@��r�";
�y���Q����6����'X���~�������Q��u�p�	�?1dXs �����C0�|Z��G���$���=��-�ַP��Ո
?�kr�X��G;�U-K}�[�Kԃ��Ѵ_���3�xK��J��X��v�u�R�:@��ZJ���lw�v�aM`ZO�t�"�l�R�{�k�p��+~fF����b�����9g>:gM^��خ(��,��{w�%\�+G�]'��.�z�%DOg?�t�kؐUѨr�ć��YX�z.���g����+�)Si}��<�^�Č��	�>��Y:�X��CR�$�N�/b���MQ�H�/�E}�����R�_<���{�q۽�u�/�D���L4{�[LM������8ģÂb�w#t\ۧ~��W�^`�޼~�ă,+�JA���S��'l���yX�&�uvfS��?��헚��H0�o3�1��J�����.~T�7��y�=��W^k	e�S�(RË��k(Z���h4/&����r<�E�=f�n���þ&�%Z@�4�υx;�u,���:"|�	�T)�iu"��W��ܮ"Eh��ͺ������n{iWp˭��8�Q�4��������N9 G����?�OU��h^p�����r~4�]Tl�/�h����d����4g�\'Ŕ�;[�m�"I.j{�m*�-�Uw��%�0@���^A�F��+!���H@$k�