XlxV64EB    270b     b70�.U)Qp�iD4pVCu�E]eg�nG��?ż�������� �]	㶆L�Z���F���N�����/Gu�ܥ^�������vn��w=�IB�J��/w��@+��^\P�"?���Y�@&��j�E���ԥ�r�7r����@P�p��\wU*ށt����:.c�[�m���= (�ݻ�ln�Ħ��ki�=uzD��٬���r����f_,t�q�n���&��%AX
F�x[����7HC�r*��!�q���Њ�2�|OƆ[T3�����/t��)x�M�p�ωH���Dh{a.�%B���N��C��ǡ��v�H�[��`Ը�� �TRX�dGI1&,T9���k`���MR�c�i��6o�oS(��k��yQ-zߝ�1s���P����!�5�+�}4�Hړ�Dq���b�]h�}��/ߠڨ��"�Ħ��tz8�7ݮzr
���X_(2����vi���z��uK�,�`���&�@��j����R����}��L���r�M'����t"��w�
 ���q,�b�<Al˸+�:�Y�*$���.qn��(�>���&}`1"�A�?��V�u��g؋a��ж�Srɒ?R������؁�kj�c�NǓ�'�+����
	�lx#���Ӣ��:¼J�-�m�{���C� �lT�<.��J�����b\���uLi� z-��xe�o����zASr�	��K�Ϣ<� �8�AS���t��g�-���+�*ԭ>��o�{�oF�����j�g���g+���y���Ӗ��Ns��g ��+�˿�Q�7.4��r���m�c��V��f�>�N�_��j������������τ_�F�p}s�a��h��r�lru�a��$m �qZS��vn��(oގ��Qh�§D�0?0R:��Xޱ�P{��J�t�E��J,�Z�\eEHQ��w���*Y��l����*���G�R���s�CW{��˔'%�oG�!?��.{� ��8�"�����EW�	�7t�_B"�mq}y��ڏg{��e��������D_��A�Ϧs���t��ܰ�x���ޚT�=�9L,w�>�6��w�8�R���VU�A��i��|�22�$���sGֈ���P�tN��.H�z��k�ZF��8w��+�*�~��C�T�]mZVP�3T�z�e4i�� '<�����
(Sg�и�B��V��휌|�%�Q��v3p�.���\�}���C��%����9a<
�b#"�C%�/pF���4�J��ռ�j��~��-P����V	ȃ#����'�-��=1��J��X25.8��cp"ꯕA���{d� �}�������C��OCUP�ci&Mp���=K�f�Y���
;,�B���5_��Q�П';Ɗ�n�!�l~<���C��
L1�q�c��^��xu�"烀..^x�)O8�5���A6����r�O	k��g��HZ�t1��؂�;�{Y���c_�&Σ��0�,��Mu�i�¨8���޺6�jH��A�7��g���c�p�
�3����
��$>&u\��j���}����'��Y~Q��%�2��+��YFRm��Mw.��/o|�j������,��h�����f�Wؽ<yj�=�Hǰ�M�෋�96G����hSt�|?�o����C��:��ȃ_`��CJT�)q����}��x������k�_�Ȗ�^�W��i�%��T��m�d�-T�N�:�x��6��j<.�~ ����Q�5B��5��I{!V�aF�(n��Qy>�ͪ7�f�N��{Gz��ԾE<������f����$�Z�x����
��~�G����0�߇�p�`���^���Gtݧi�ZU'��``�`)�ˑ9�P�f|���V�Ҫ&�I�4r�_��Z
|����Q�$7�W�z�>ll����ՠ����w<��s�$�V993�vC�g%Un���t ��Z����hT�b:õ���[ΩD7G�!���f��U��l�A!/ ���AVd5k@�F�F�FT$�o���ȋYy>}�����IN�X���li�)% ?^Vw�o�h�q��;)9���f��ǃ��٫�P�A�%h��X��1�Fu��*S=�V��!1x
ڨ@�ҥ���G�j��P�ћ����wǃO��hΫ�5�I�,�1�2�|Ok�������=�r �r��|3ѿ�����Uc��S�ҋvsJ���*�6w#'���z�	�������#�[��̧��o���X_��Btȣ���ql&�}J�ʝY
G� a�D� �÷XN�Wrc��XfS��8���]���W�B�,s���&~hwߺ	��@DW,{�$�򊗔�*��NUC�L�m]����
�	�K%Rh����dχ�A�u���M}��3G��?7�`��,L��)���c�O��5R�6�cU���s_o6�ݕߛBL\xB���C�j��Aҙ�6H�v�7�g*�<�K�R�c2����`���r���,m�����	�7{�V,�:��6w�C�j���=�`a����l���A�����G���>��W[g^Y�z�n ����$��F��%�q�O9�+΢; �`a� GX?Ѭ��<z���3h�b�N��1�Q&{�GO��n���!�� �&Lz�P3?۱�Ez�B�"eyw�Q�z:���60I:1�qs�m֧s��!85����ei��x�$��
�e�ժq��ԡs��>�}P!5�2�a'ۑEFh�����Yߧ�{v+`
�����ؒ�;�ʚ�#��q�� G\ 0������cQ��:%�uN�����<����v�!4�