XlxV64EB    2e86     cc0��:�܌�G���o���_1���M����ON���!��监�%*+r&����q%���3��_��_8@���#�Ӓ#��3r�U�"n�����A�O�,�E��pa�Ys����aߝ� ����mUm��}s��+.slO�ϴ���6qt�t����-񥏝m-�VtNFq~5'f���}�m�����"v��e�B�	x��wdT��������y䎥���uj��=�D�Xp/y<[�Ky�� Z�Uz�{�d2�t����.��ހ<�uc�+^h�ҍXi� ��Rv�z�a�8^�t�`'��Vd�*8�Ř��d�A�3o&
gXC���~���J	��+���d����t�2��xC@B*8�]pM�����_@Lw-�^&�r��C�7ۢ,���M���:t�b�CÄʭ��\~斺���|s.V	p&7����a��p{2��dcI�,��;��a#�}���È��K�_4���^�����m�K�9���kZ�T������ܝ}���lĬ�X �U��U���I��%�f��@��$���	�9!�[}��f�o���^CbҷNծ�����+_�:��i�����rb�U���e�)�H6��Mf (-��8 XB�Y#����k�!P�����<j�.e?�(�~
�R�����&76�S�J��˝��?�ðK��C��kV)�?��J��{9΢<�!GCb�F'�c%�sk���!G P̥rf]I'[�R�U��t��X�<{���]c0�fI�tړ��)l�(�/����֡�<GuCl���4:~E�hH¨	�G`��%�j�@*�#/d���b�u1�;�7��E��g.X��|1R���/�i��%�"߈�=~���Յ�gd��uAճ
�|p��C�x���8�0���,&Nj&0_j�����/��p����g��ˍ6[���x7����v�̅F�_kx�VC���w�r�qا!����	P��Xc�$�1�'_�i߽�I�դwN߁�w�k��kf��Q����B۱�t5�E2t��}�4�f��9���J�8�6�"�����L��s��H!��-.�L�:�W-#���DC�����~`��V1=����p�"_*4|�Hj=J��L���$�9=C)���F%�cjU%��j��F��fx�R�;� ګ��*���nF�䵶��'��0�llkp_�=��M��7�/�4�[n����Qݮ|���Kxj�H\B�������ʷ�\R�e�I���1��H���_��=����t&�]�� �x�H�a�y��������T�GBZ���J<I�)<Hņ⢈p�L�X*6�9!Q�@����Y��c!5����J��L�x6�	�H���RkR�Kѐ��|�����X]���9�v8sp�>��\�t�an:̻�S~��Ht��3�7C,-�3�bK9*OW
��T����F��+����j}�{����T�$�ެ�9�n[�22�����Z4��I��U21�+)0}ۻ��Խ�SW��jP����V��3�/9�`ƹ�Q�8�K=j4n��ۿCU�hĝf���
6��%��%��l�Z�ߖ[B��>��>�,�ft�8Q*�|����+vb��4��sӺ4��*��ĉ���:�R���'a���}�_n(����S�ɬ��gq DV2Q��h��8�;�̫\��ڎ�-�;�1������k1��B;f=$}	}����z�u�͖e/�����6�%`
���%J�}�x�#y���Y��a�I����ʬk�s�C�����+���
�<D�o%-!�8pH�����a������2�v�!��]]9�6�r9�m��`����S_�D?�o�6���z]��E��(���%�b��zՄRړ8V}coX��R��Ģ���z�&8�ꎑ�=��O6w�<�s;���7KK�V�V<N���|$�3)��{��̭o����`&��*&�Y6�}{��ZkU3D�7��\��%sRG�w3�|��j5%_�#�)O����v����p�f�r�^��}��J�.��h� ��z�+<[)װ��Eіl�m�����F�r	 b��$���}�j��[��4V��j����#�?(����>r�����4��"J���fA�ٌW݇U5�IwGܷ>�cI,�ӫ��\'�g=�Y&�C�pkM5��|r�~Ao�y(v.�&��Ii9HЈ�⺲q�H��͖���
0�u*�ԩJ����hU��ʹ�����N��Z�k��̍àpjH��<wV��Y����B���t��~�tw�'������J�z�ې�#N3sѭ����E�٫��J����Yx�]I�ŷ?���5}D��&;�
�Fd��LM�	ǳ��t?�F�٦���K�s�1���WX����!�Zhg:���f�e���A+�n���L�GEf\u@�ץ�%'�m#s{i�9��+�����o>}����P����ok�Ncg̕�[�`X��H�T�Ȑ�9�OS���7�`ݐf�=Dp�,na�L�1���:���O�1Zb�&9]��0	 g(�`9R�lb�[ViIu����*��ݸ?}��Ή�2G�4�=ć�o��E�:=_j���)�y��'Q��װ��R�J��ULe+�`�E�*,��Zێ`�bx*���Gf�(2c&�w,�r��$�̗"�	8�N�:��p�	�1DS�5��,r�.�ǫ|�	���~��#� > *��;�t7�;����n�t�\�}X'��,���~(i�@O�`v+�=��T�����'+�Y�s<p�W����;w�7�&�X�ӕ�7��jʉvlm��4�j�H�:ʀ:`V�/�Q4	��Y��b�W����q��0i��C�Z�2>��$������ũ�U,��{%�b!�o���¹A���V�;�[m`]4��o3Y&z�g���X(j�z(�h�?L��Si!�7�~���od���B��b��9�>k%x׏�F���S˧�3���1��.'5��g�C\ܙ�����6T�f{�e����;bޖ�x�Vz�M�05�
8���i��9;6�Y���^K7����aQH�ɬ��e���'�_��5[ph9%.]�P�\k�^�B�-'���<;c
@�FB9�0U��̀X�G����
$���n.d�d`�D�}��a`j�n�ט"�9��m��\��noR�0�&