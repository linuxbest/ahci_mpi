XlxV64EB    15d1     810����KD��]e�Yf�����/���7Λ~��w 8<�>�BZ�-�E����#B]����Y��^&��7�q k_h���h�w�{i����[��;��}{*��z�4�ܸ��v���۔>W��»	K�"�Z������}g�@���*�տ�e0t�L���(_��M�/`�C9����Ă��i�]d��h�*�}��mՈ����BN�O�j$�wU׵�	��{��6�}t��d��o�v�W�i�~囥��@�v�(�b�>��4�����k���2���T��B ���_ ��T��_��|;eeKHJ8t����ܝᓗ����j�Bf��2��Q�&�����Z�?)���lGx�!��7p�}Dd���E�a�z�n��ss��*����h���v-��$A`|��Êca�|Cbfa�¼�\Ax����i��"ȅ�̌\�S�#G�3��:
�ú��ţ��fQ�2���9�	g�L�Q��fJ����3e��͈�_�I��3�xylr/��%N��\��+��"өN��I���4�_1����%S=ͩ�h8�ѝ#D#G���M�D ύ�`0������d����3�Ď���殐1��`XxJ(2���a�j���#����@��o�|�c��g�=���u���}�gA�s@ګXk�M���'���	lr�k3��6�R���:���ʢ��뫤ӯ.��#S��H�1�+dpf,�ێ��L�U����0��!\�ڥ�&#��J[Ͳ�w�?�6������;dZ��UE(��[ل(y������V�]��'^���5c������H ֽ_�2r���fB�0IL������T���Lxi�tT(��w�߃�qw�	34d�����'8W�ޏu��H���FA��}Pi���o�g�zhA�
����n�W?#�4�9���������]��Q��=$�r b�����;�vv��L��(^�_VQi�I�-SdQ~�Vy�g�N-<ܤA8F+��S�����͎){�Һ:[ѢuӀ�>f�Nr�v�q�7/Wj��m�B.��W!�d,#1�p��ч �_K:7*��]*�|ʑ�0�&����>�Ǵ��Ej7�~Si��LJ��Al�6mW�&�W�9hN+�wdfJ�X�O簫��2�g��)��2�������Jh�N%��!�aX�d|膑��?~B{����G��H��v�^l���B�p�7jӍ�vO��_a��R�c�sqk�;b�{6f,;�F/�ݻ!F-�.��6M�p�*ڵV�g�3�CjC�u����[�CӅ@쭷�X�{��(O�U��X}|�5�f'����^L>�K�z&��C@-%���$�ÜЦ̑A�X�2��K$���+h�l-�3N���] ܮ�+�V)�ߗo��`)�i`&5��j�2
^N�9ή���{�O�Hi�"�t�A��KҴ�^��ޘq!|�Dch����=�ެ��Rl��Ʌ�������l��ͬ�N�[EŮv�l�<����'��V�hY��X�<(�I:��`��T�U��T����p��f����*>x[��	od.\˹�G�ɦ��+d �H�1��I��tA�:4S�K�*��Ulw;@����]ǿ�7�n�S`Z^ǹ�ΣT��A1���X��Y^�"q���0wG^�ԗ0�
�.�!l�D�ǋ��],��
�~��W�uY/�,�^�5�4[���@�w��'~>�����|�\0����g�Թ�r���ȿ�4'Y�4�,��.9���@�=Ñ� %��k�g|�����:Ou�i�ʻI�?-)�3F�Ѫ��S�l�����D_�~��I��U�2Z�!}�׸G�������r"w��[D�h���
����]�Ǟ���v �����}�O���6��Z5]��h�";�#��b���	V13�M���+�K8Ľ�!.��${���LH�f�a�d�2}�FM<0w���B���{1u���pV��7�S�
�R#���tF�g��K��J�\�1Ͻ�Fl/i�e��2ع.�l��<