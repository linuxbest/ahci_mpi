XlxV64EB    1fe4     9d0�T��aD�b�i�6�eh��@�>�X|���:u�i[;���l&|�@]��o�6F��>��o��������Aqf5 �M��q�
���~$�����ceR|���[�S�<)n�=Ǵ��,��J��(�Jvʛӄ�ٹq�S��1X�#pi��ԸG1l��4]� @�9-�-s��},�e&�4	��ͫ�@ز�!��>L�mmYox��J?��
���lzip�+F��P�џNv
b� _' ��p���={��<N�e�Az��7^򵱼$B�H[�.U?�92)��Tm�B�qoq�|�g�)@�t]*գ6e0X�!{w��A�P�A�T��-�>��n
���d�4p�5�T�Ͻ��}9RR?�CGU3HQԡ6�z����z5��f>�pa��K�O��������Hv�����֡]��ak��t�'�[�5�  ]�p�<@�ʓ+�+
�#�h��'s����
!CY�7�����04�S��rj��򈊃>wql�w��1w7h���E�����39l܉�N��3����d�P��*��{7`zm�Y?catXb_9�Yr���r.D�t�z� �if��5�ɩ"!�8�WYKй�U���[���sA{N#��� ݞ�;ug�$эx�s2Ѽ��B�U��>�n�AX�M�~z�3N����y�)o��]�	��eN��A� 3*3&q��ښC�氦��٧v�OG�q�
CpS�a7��A���l�������A@�;�s)���'�{�Qf�^�EQ|�$�*�����K}{��$�a���o��/
vv�lx��B�H@"���͚������k��B�)�Ħ�ד:����q@��,)��bѤRE�G_��=�\��~*t@�z�e���]Ei�g��^
(����*͞�i"����A�6��mB�Dw�@�X�_�2CF>�o'��qgO���k��5R��%j��]�������i$��9����{��'}��0��s�)��?�����'ՈD,����د����}F�Ȼ�|�2]��n��ʦݒ]���`��cp�"������};��R�C�[���<d.� l��:���C@_h~|󍨙D\������S�<�sf`p7ݸwf���
��!*�R���@?Z	��L����$�����1�Өü��p�3U,�\ف��ں��"�������c����ag{��攠�[�=�b�p��a�iL5�0�D�D��QM��=����rxy`�:�%���+�#7ۉ<8��e"����S��x��=N
���9�0��;c�T1&lK��$<T���m��>
a���:��I�K�.?��;�oW8�Ơ��dKC<1^^~!]�@@+��w��N�l�=d
k:� f)�P6�y���#��؈�x�x���Y���>/#�
�ԍ�"�L{�M9���(gv��|�sM���[ ]n,lk��͔r�8������;� ��0�w`�"i���$�ޞ
��?r�.���ǁ���4����
���`�F������<��5�jJ�$51 �en��'@��ʬ5Z����"�	�TO����G2&o��XQ��g�V��$���R׍����
=�a�jH8osTCL�`��-�OW*�����r�pNO_����O�lk�*b�#q�nt����P2���:�D�{�B�����;�8F઱6%p�0�Į���sM�e�6�
TX}ۑ�/F�����D�-�~�xc����(#���LҸ���PH������ۉK��t�?/�I��<���qJu��?��q�||JZo1;EX�:��z~J�4�7` (X��:sF��ցu��I�?9˳l���� l͇�]U�k��P��%uŢ| �Dvn���R�Djí�nW,�{�a�'���M���p��J�Y��dg�����#n6���ⴋT��:-9�c���[�wT(��XM6�����.k������h���Ds�j:ʯж�s����E�~X�����v�U��C�alTV����Sz��.�f�+|��s��T��^0/�eP��~p⋝3h��
�)��Qx���b��:U?�5�0��J��Vя�Z%Ǐ�U�#�ȃf�><�ز�H�݋�ŏ��-?��]��mC|�6�������%<�i���(�&cN��k�H�!��$�Md�
�E�{��9Y�Ќ���+�ӹ~�EE�iB>Rx�7������X�fb{>Q&�>ԫ����>�S��_a�ٮ;,���u�.�Cq��>'xg�C^��]���$�Ū|I����P�1�9������j�B��X�u���Q�TNjzǲ�u�tBc�:��������38V3��*ۏ#Qo������A��p��7�^�?��%���?Cl�3��ְ��ӭӲtU*rĲN ʅ���"�iz�߲Rb�>�k\k�Ȕ�)���I�X�b̵��*"�b^���g�ۊ'�5*~Č�/�>�\-i+(���t��:��F