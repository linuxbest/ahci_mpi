XlxV64EB    26e0     c00�'Øy�,���GG�o��:�DѽSf�H���A�,U��)�T��ynF�������CE�h�"	@'0P��u��j-;v��[�RJ��[`>���ޣyϵ�Et�ﻹ��C���`�wx�.�@@���{J��s���3�k5l>$.��'䫷ٿ����F���+����Qz���|��
��T�_�c;�73�lY)�2�0��S�� �t�T�r�a�W��o��E+�F�&��F"#F�(B��0,��_�}���N��q��x
7����*�ͼn��$�噀y0��r�|�@� _����aJɰ��i_�zb�/��{��R��u<5�'����<�:��m�ḿ}�!0F��Z(���DUq�>���c�A��s��|��rP
������:��@��|�O��Y����}1M�Pnza��:=�=�ٍW`P��E9���D�x�?H�w6�sr��k��0�����ģt�3�j�B�$e����-C�3��q�{3yU�FN�CVLc:����ٰUj.�5�-+Z_OVB��F�ĊJc]"�q�W�,jF���s�:h������0;b�����zT���PV.�]�?���a�%�ik'����Z"�v�U��@�k�4t`�5���[�w�^��`����d�p�6���?&
늋; ]�H�MwF'�NX2�D1�=�f S��,�I�i��liʅpv��M9�h��އ��s4���xw�-`��ۘq�)��d�_F�n���鯰���ð���mU�0���&�B=.�"&�	��ݔ���Rqqt�k�=��e9�S���ԝ{F�E:���؝ܚ������3�7M�?C�MVM��3��F�ܗ�}+N��K��i�ޣ�Gt���M��,G��}�"L��}G*۬#�v��_�s�%ɻ'��(,��Dgrݩ�E#HX��O	^Q�72֦�pұ��~��٭��Е�óN����[g,�-�@���+�ьMwe;��O��`#�3@o�v�: �S���ؿ\�v��������_�E�I{#/�JLH����T��~�
n�fx���,q?� 	� =����#�O���#�FV�l�_�{���׼J:H��U�AM��/9�X�h����ba���̱�"^��fmkء��|�wq��	�J�����Z�� b�S;	�q �b`��]�F��l�t@��~:�ij*�����2�z���h ��f톁뿽M�vg�ҏ?�8�T3��F������
 s��<]'���(gk�"�I�nM�n����{�}du10!Eo@E6u&̾I���p���I�k���>5Qw��<(�o�d�r�������෴F�7�:Kn�5�O� N��8вA��h��PI��i�"���%�A��*�p�3)3�Qq���P�m��ZǩoJ�;�txq֧�tC����?9uM
Y#	m�!�V�������<�M(o$�jd_�u���D��ňv
�@��<�&���1f�� ���f����/�~>3�����\ �=���⧬�F��J��}��
���8����0��č;y�TE��T�ȅg?�����t�+c���r��4{���I�����7����$��"p�p���q�sR� ��/o��9���x��e�ų?�g~+�.�݇]���;��(���1�(��޳C͵j�FH���v�,g�D�0��|�|=��(��yt(ڭ�|������	��=�ܘ�b�+P:j	�G9x��XQ�Ȩ��4��O+
�P�x_'3}�[iMD9k�BJ`�7<��a�P���s�\^ �}�F��;t\����ꎷ�6�bO�����;�臧U��Q�%�b�� �-"������%O�੉�:bK>dd��_L�uE�A��D�Lxr�����C��5w󆔄���e}���7���[T�1����u��̀�G�ȾiJa��i�ΓS���.  .F��&���`��)�z�u���<t𿂄0�ҩ���� �S������Ҝ*��J��"bd���*��MMɱ/ֻ�����(�=�	�X���ZP$�40���6����I��9(�6j��)�s|/�՝~]�A�_�>�(�)�#��'@(�[��`�J�	��k�aN�z-[=|w��䶫����|9r�mȷw,Y:�f�#��غ4r����}�* �N�#��?L,4�k�P�B�w�d�9G�Cd�ƞ��/ � ����vl�$��R`�ā�O#��Pb�M�ƾ}��gp��d�n�Q�mѧ�&��!����֑����kLn�H�kN�y �7� 
\�#���v�+�J��}P������Z�2�� C���{1El�r軁n] 7�-í@�H~��X ������z�Gov���ۙ�O����y�f��=�F��Z��'��ddFm
�9���H�RR�o�YW���B�p瓪g�JIO�p����7֝��N�JzV��5�9��;N�PA�ǵ�w~Ȇq՝��}am��o���L�©Hϕ�;�2!�aFFIL�拄0-D��s�(ϟ��t`=�~1tzq,o���l��4M�Qp����h���58���^����e6&@I˸�5�� �H��-��(�gܣ"iWdN��{v1U[_���m�� �M!�M��ɉNpb@27���\���c�=0�,�jTT[�\����ۆ���*e���*��Oc�v���t������R)��^�j@��v��;�4��رj}����'�#G<��}�o	a^�t�ޫݯUvFs'�E9ƇZ��	�ְ����1���d��J�LJ"l#1uت-��/����]C�~��d=uŇ=>�Xw�ɽ���Yi�ѹK�o֨�<�gs��D��B<J�e9�#��f�@݀=���#�W�coۃ����x�x8���%9�<�J.��eu>l���>�&���q
��m��@�/M�dd_�$��:Rǉ�~�S��->n(��]jŭ824�צ�h̅��