XlxV64EB    53e2    1130<�͡_�����I4H&
V`d�oW����#��j�y�,���4C�(�mU,�`L�� #f�
;�՘,�5���_���r:���������@��9���5�(!�=t�Z����+���6UեN_6Q��\��{�\}�]7�<6�%.�\Q3T�w�Uu���7<(:��+?9���i�C�=Ye��xG������g�7ꂥ^��(�lڗ�%��{�hO�ҋA�MAL0���i6-T�ݫSlz�H���	�w���I�+�|OO�3|��b�R{R���ER:�;U,8����G
�>oЈ_K�L�R�	j�6#�VZ(�ޜ���:~X�������Fyl��nH��Y�y���x��8���^�
��2�Kл�����^�J�l�п�n��r�Aw�&V!��
�횊�8-.su�@���W�e� ,m� �q���8�� 	n�L���(:h�-�a�-,(����gL��a��]�"
��>I�'wܑ�*�RXi�cM԰{BK$������ IF�$����Z=&�3�K�����8�TXO��3�yVik.�&.�1�Ê���D.�Ȋ�f��5q)Q��=w�����a!������Ú��8�$4=�/���,�LA��b��V��b�qY�w�#�s����|$�Q����DZ��ʌ#��n_{(�퓚c�*�oO�����@�"�I����]�1�:�y~
װ��o1�[Q������4M�b��斢�*ya��	�TY��S��Ά����D�;(� ;�ۉ�⤀����T7�h*h�hz�ކ��$�2�����_ �6�?৅�qe%X����i�� �ż#�4�*\���Z:
X�U
��z�:����:�H�Q�%���2�4z��0�Uv�C��-�]�HJ#�c��A*!6=�Q�֛VE���K-�A��`HS���}�N%���4�~Ȍ��g�a@lGK<=x���&�3�V�~�o�5��|8���d��kAvl�5Y|��O垎x��<��:�dn��f�YV,y��E}����ʤ&���h^�bـ�-��S ��*Rl� 0i+�ymZ��쯕�L�K�ХB�9�8ҥ2��(�k�G���Ӈޚ&�S���ё� ��[��]�;�o	Eey�٤�`U���5)����<lETÈU5C�''�Y�w�i�4P���0��飵Җ�(V��t1�7�o��?$I�("�x�d6����CD+FBO�e09��� r������Ԏ)��*���xO9ˍ�ΉY��[Ɖ~������M�������{�_����&r]l���1?S~.V��CsbkǊ�(7YV~�����,o��
 ���p�m�K��8ؕ��WA��"�9���z��-Woi>��1�Ýy�V����a&׼���9J�k�<���q������{���OH�^�8�bhh���騴S��x{�g��Yr��&'�q�p`��ؓ�����q~��7�e� �{�k��Er�*x�`�}�R�3`I�j�ϯb���$)5s�J,s`�cr�u�b2%8z4��2�:��F�{������r�j�7x�́�����n$W��6�X����jZ��˜��Fd>�%�P؟��d��t�ɵN�Ó��'Q�+�9��9gqL���&P�RxG���J�ͳ1l�ݖ4h�P�O��B�'��5�;�+x4ܾ�v��d����z��;:�O�E��>x����6�#��V�I��]/J���e���#��q8Z�>�#�;��$x�豣��5.O�<���4z#։ʷ���v]��y���6A��x������m�P0Dv�<<u�eq�x�<��[@�H�"h�|Y�f��t����
&�9ĉz+��l����I��-�ޯ�׍3!�H�F���7w����s��Z��q��x+�"����%��u��ix������6���	q����}V�#Zv��mV���o�AyW"޹ n��{��w�Tk����(:���[X0���`tU�aαH���~7G�3����!m��
��a�-'�I�;\���޼�92�V���y��s��V�@���*i[	aˢzL i�y�����id#DB�YF�>�,��M4B�g^%޲��3M���6,��:�e�4}
e�{�dYV��1�� e��&��9�mN������������¢K Jɮ����
W���!��M�1�?����%�u݅F1��`��H�̇�&�2��j���:��P�����e�K|=�f�&+H��.)ԨS�D��ɒ�glѫ\l�$�$�,�~"&+%��k:�3?l�U�J^$�$wRPXѓ��\�������JGx��k�Ρ a�	'�t�����C��<9R��$~3'�
5x���v3-�&q>]j)/��<�c��s�Cm��*n��KH��l|�?y�'Ҿ��K�['�͍l���u�*���2��A!OF_i��j������Y�i^��u��/�68^�� l\uq�H�_P��7�wk�f�ߝ]������P�3��m��,Y?8���8���[�[Gщ��y�%��K؁	KȚ�R����U�K�O�YH?2���.�1��LfC����;�IĚ���&`D�� ��F?pԔh<Q� �����)�]�2E����q�|dy�3 E�SՅK)�3\�N��}�L7�xo9�`��fTs�XNy3���JWpNB'F�3�:B�%�;�u��]:��E�f<�q<"�2т돜��ǗU'��_F�+����y��X�M�:
0�Ҧ�����O��Nd����[�W�<���w�WU��}Ca��e���T�3'W@F %Zb����SW��E�kv��b�jaPՒ�o��'$\��n�Ћ�nS�]��ٳ �(r��m���ɂ7x��~��UG�0]+�ٮ,5!w�"{h�lh�c�4`���J�u���� �oW�2�S{�n��V���yբ��/�^Jp��=}7%�O2M��W��c�V`P��"X(	F��EW��X�qU5��9D�Y�Y�3o'4����i�jz�l�3�r��"�T���$�j��s��R�H�A,|S���fP(��*%�ؚZ��]���w�ұ?:ڟM[⾑�=6�ǪZ�;gؑ-X�<^���[z�؅7��UȅEa{�����I����?$췤�*���U�k� ^M����~Wo�C:8vn��� P�L{+�ā�M�j�
��G��yأ������y���+���ƌ�E�(�q�<���N���g���'������:�t�O�� �u�ܬ����m߽�ue+ �j�S����,����|br�7�9������y��Q��tuE����𽃗�7�^+�oG�^���~�(o��$D�G��a��M�^�ږ+Ga�5EK�FR��=*QmJb��nr�5��*3!�5�l��Mi�F�Xu�r	�W�߫�*��6Zks���@J9ah�R�]��b��VAM��OZ���Zy;���qa��<�������e����`ەi�Q�o��gN_����Κo��M����ء�?cBH�/u-K�x�	�Z���޶q� 9V�������O|'��3WO'��D�R#$�������(���Iw��u�=X���S?�Ҩ㲡� �-�����Z���9��*���Q�P��%��*�� �>>�kd÷�ͭ����4\?QҳNNԝ1q�? e!P��nY����/�`)?�(�-��R	2��<�N�*���-9QN|=/��q����9��&�:�)�Թ�O����S4�x�B����j�U�i<��[��愈��U�S��!	�Zx��wv覴(i:��S5ɓs?0����!���!gg��5�=���]�"��Yv���7oKr�l_d@���M��a�&��d	S�jc¯t���Mė9���oi������m��p�,���"��ɵ���0��~��i�����p t�O�XGP��[�'ب�{���rY�����
N�kO �ų�ؐz�!Xa9L%�C.6*��W�_�*�mlk���>�U���`��N�A,�Lǳ��wـ�z�@���Jw�^�>����ĔO�>M(�5P�$Q��I�A<�eԜW�0����H�c�\_*(�z V��B���:�6l� ym��ODR\5����4O7�~T��t�ǥn��-÷%5��5�Ao,5Q������m�!��W{(�mSs��'�6���8g��{�@օy1+�
P�I_�g0���e��Id��(�s?�����B3n�[�rOA������k?1�[�-�ݲ(t