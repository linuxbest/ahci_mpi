XlxV64EB    3366     cf0�T(X<ӣ���J@����0����P����*�DF��h7�&ǝ��)��g�XVAa/NKx�l>��@��}H�u:�i�S��zp 󻏑�o��=� ���"�F�2�J阧�ˬK���
�3��	t��w��W�DI)Uwu<b�a��m�BZ� 6��D�@��ұ;z`D�:�Yx��Ic0j�ל������m�w ��dq�=���* ���?���|�x�:�䌙���b>k(�`hG�?�q�Gm+�� E��9ק���VB!��v3�cY��o?�:m���8G����u�0-�C�`�t\\O�������c�
A���Ɩd��*�Rx�eQ���~��L�{8����w�?�?�	��}�$c�����F��h2�Ϧt��<�R��~	�5�,Ъ�(��u��R#}��i�Bh�&��M���z�X~)�����9Z1�+]y{��i륰�HX|ߨu���aý=Np�!<K�)��L��^�HzZƝ�ga?�(GW���jj[�e��-+j&����3�x��»LG+��E�k0�;�ߨ~-�~%���ҥ�?��U*/�ͳ����~�%�&F��]+����*��
;��m��$y=�/	��4�6/���³(������oP!�ķ8���S�1v�_ȦT#��G9����"o=�0��t�+�0ڽ�REPx�g'krt�	����_�1�c
�^⏺k��{;J1N��Z/�2+��´%��=��r$*o�x�<���2��ŋx�Nq����Sz΁����;Λ��N�Z
^�!��x��D�q��T6�WV��yP�p��S*u�G���5�<�zLa�TŒW��V𤷃 +]��d_ z�H����cf�;�p,D���@��;{�k�""C;�N����=O�a�X����fm��@�[���4�� fm��������|��Vd{�H ����{R	�����{b�]w�.ܚqY
��^��GR3�҉k5t�:Q6*�G��kW�Li���o�J��j����<j��,��K?������~��J=	#B�u�������p�9�E��+�>\ע�ٶ(E�H2j�J`��Ka���OF,��R!�?�:��[�<Q�o����Py]I�	�$QM;f�ǐ����3iݶ�j��)�x�Py���k������h?F�hRa�b@mD��8���Ũ�����dbA�a���BC����Ǹ2��]ԩX��}ų���,.�A^��L3;�%��8���l:�����łS�	d����%��L��p��"���fP&M��K�����N����m�C;��Nte�}�Ҿ��'� u��4��x%�N7@��مA3����ep���T��"�ۃU�i�Ksǧ�-�>��E�� o�,�$�A^X��L�(�kZfO�0�W��<�-~���������8�����瞹:s�5��n^��;7Q�W>�<=w�N��J��S9nF�����K(Xh�Է����Q�7�tH�� G;��Q�Oݗ�DDk�V�L/�rl��Q->�2_Y�t�i��d��o���������0�����`m���S�m
����'�ZZ16}�]P:��5�n1��\��ɵ�J	�(q�0�2!�����l~&�:"�I��]��km��-�N8�ܮY�h^|!��I���pJ9;�ճ,��'L2o�9K,�s04��-u�f���ߩ$,Vۇk��S����Z�-;=$wF�Z��]���Ex��	 �c9�z�����)��Q�kKkI�vCls��[{
 �~O�	��0��'�-��J�P�^Y`[���_�<1�GfEܾ�}�+��7Y	��Ζp�޴"��~gz�����D�GW��,+���"_;�;�es� ��HF�ZidB/Z+���3Bc�cȜ:�7sL�&�����{K�ǫ5��I�0� ��$x#
�RX��`� b��E�����	��J:�g�V:���'�O: �V��W������'�W�8YB�3!�:�:R��C��f����0��S����t�)&�/��/U��fuV�V�Wv�>G �Q.Φ����@����ȅ�g���B��3�k��LC~Q|1 �py�5��E�0M��?�^��.9��~�����X��V<5�ARr0���G{^�d:-3L{dM��0��4��tw��m��9���������J������S���l�E8��w�3^kBx~���9[l�q������96��n"~e��`���)�Gy��Rt)���i_����>>��aG�9&t��t�R�M�^їᄛH�	�5��.�Ki��P���k=����p�0�?B�M�i��o+��wr���P�[QҴH��K%л�Y�u�܌!OVe�O���!l�ĪM�x+:�d�KBЮ"���ٲ#'ǯ^���L[p<v`j�2�	�TM�L=�*[ʢE�k���*82�r���{��,�w�JU���}r�a�4����p&j)9r���^1�� ]��/7��q���--J#��b�w��Vkc������`�2���]��]p?1w����Zö��m>y�����.��������n$ŝ�4���I¾z����:�2*n>)�S��r�R��O�4=���~���\���1�˯�4A���4mZ
��j���&c�KD}�N���WN���~"�Tq�xVxp��G��$nz�Py�!+zO:�7��
}Fګ (.n�x1h��7M��3?<�O�_���g��D��?^LU�y��������'D�a���d����zN��qQ�0�#Q;M���ô�?������J��/@y�͚��UCh&����ȭ`�u�̨�9�/ح��d�\��P?�
�|�qX�\t��9d�L�Z�5�7�H8Vߛ��@��O�,���*m[����v��0'���z2��H(,����E3F���S���H���XX�I@* =j9��s�w:�b�}G��Rl�����MQd��6~P2,��bcĒȻ���Ao���%�\j���2|�p3�V<��H��ͤWf�hP@ׅrze��t�ZcבNjف^�F9�k����R�����h���F�H�{BR�|7x��,��/|Ge��7Z��I;�wűC���x#�F�路t���"�q���� #������k��(�M�sIX�g_βؙ$/Z��d^t��ؔ�;C�ڮc�G��x����ȱ��m�*9?��#J�'��j�FuCd5�q��B|���K_�Jw�>e%�E§}��� �-İ��춰A�9����l{_��v