XlxV64EB    1870     6702svX�u)F�>�E����Uo��*�q��y��p�.A�fVU����cϧh�'��{�M��	.�ޠ���z�3��¦��/^|���K\�l���Ԇ"F֘�V�����H'�@���bJ�5�r0��⼠����A+��r��x���"���,���e�P��sQe�w
�_�{�::2��jnUt��Ny��ܾ�z��o
�3��W�o�<�R}B@7{�)U��E�q����V�h���ƹ��T;/��32�v*��3ia=ߠ��wu��g.�̌�9��r���b�f�y�07!� 1��6G��;2�b����|��g���rդ�DyY�xU;Yb4��Y�u�"p�(�N�`a4'�:�Z(��@v��ZO)���#�U�)A)r����hQ/\/�>6�ݙ\b�o�iF���G��."�=O�}��ؿ��4�'��f�CFہ���g��M"B����L���^H�0�t�7�eҦ���`�8ؠ�)�0M�V�S���J��$7 ��r �*8*�D��@|��C����X�x�HwT�'@F���B��')���J��Y4=������+�CU�~)���D�Q�:��0���=SC�i�� ΝMux�>���B���������䞌�U��!@�`�	����Ҳ���߉��F7Ht�m���q:�����[�+7j��cz�z�E�������Ŭ��Y���u�3鴠p�	E��4�U�d<�p��;f�7��\��D�C���߳��^(���wk���rWc���b�*�a��bk��n~/�n��7�����"�Y6(����>6s[�s&��-�Vx�P��Mڿ�7�^D��<w�_FI��#	�+��u)\FW���y�<���Q%m�N��Y�F6�1�-�0�YO > �ĵ�{	������:�0��E>)n��)Tr64�ɖ�h�4��?T���f>+��a�Dlw�U�d����N����G�����:H��3ih���]�:=
���tb�k���ܶ�5��D;^�籝�H�Ü���2Ѷ1��/"+���b���#֧E:YּyYKT��BA��V�@�vB��
?���D�}ܡTT��E�ϩ�+���I^j���z���w9$�����?q�0����4q��K�/W04gz����Hh�G~i"q9j�I����Ɣ��M��i���Rr����A��.�9��a�̪M|6XQ�XӔ���T琅Z�>��}�I1��!�&g�E�D�8����J�|�4ù<�I�`�� �o�W�/	Sp�,=��LD���/��'��Y4j�w�⅑���8�)Z�<�2z�16G�=�āAV�/~�sSb��i���yH�Qwgށ�����?(TQ�T�����n�ҽ"�l�5f =�[�[g�`>=�7-�>�?aG����h���ֹ 6����n���w�H��0���!~�V���B1!� s뽫�x*���j�~���h�9�ySL)о�/	Sr�����I}}���$z��,찲��? ��sӤ(P^=��cj�:̘������5u���=��k�
,�ȧ���㚠C��V4br�v������&C-g.��rS