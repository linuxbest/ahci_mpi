XlxV64EB    fa00    2de0I���~y0���(ZVE�S������!k��7��h�D�^�����G���-0�J�n����B���7�g�e��	3��B
�AUtEff�0l��t��������6�eLY#�35���Sj�NK�h֔�4"l�K3?��j{�K�%,�$�<�o�tn��-:�kh�'��-qx�ҫ�@�����T+���[��N�j9��] =�\��t��w�wr�矩�IȥW5}D��gX�T�J��<��\ݭp��f6�CX�V������m�8{�L��c��,ꂱr	� �*���C{)sێe��2���8T��6������a� +��1��#u�t�&�0��Օr�ұ�rX����t���~YO/����:6������}�$r}qB+c�T�IlK/[� B	�����>\L�<�J�(�y�Lg�]���owW��PE�O�|�˽.���U* o �qjGd�\eg������CA.0�H�贴���:"��]M��
�)��Af0P�Nw�;�
%C�51r$�u�:5Ё����x�H�0ƤC��b\m����Z�c������=V̋�q�k���PN�'���`����T��<�}A��F'�E�v��=���E��!Q���"�/�L��@a���Df5�:��'p*F��$!�F�۰���`�&���ryl� ����L�O�<�p�+�}��F�ڲ������x�$m��L`��۾�.T.���Z0؞4�JD>�*FG ��H�l�.wq���Ņ�*����%�W�����rb�x#c�Hg�4%���`3�cw����k\YD�q����� n���^Eu���n��1�p;F�ü�|�v��i�j���hzG�F:�ˑ��@/	̋Υ>PO"8h[����OA�d����O�Z��o�T;'6N�N^����[�USֺI��i`-Q`S�J�	\,��٩�G&������	�`���{�U����Is̥�9[b䞮쥕^�UF ��c�b�t���<�'h	���:�q�E�Hjl�ֱYu�.5� c�Lq�'���/Da%]��r�v����(�h�_�k�C#V�=O�w�U�{-�2�+F�t�J��d��cV�׻������_H��T�9�6uT�nR-�'�+	� q"������tIr�s��Fc�l!&��F睐.}A��7�`�Lk����[^�����<��(]��۷&�� �b=�y�̪X���������u⫗D��f��J�jV�����4b��B�$@�Rp���,���Gc�i���,��6�>2r�d���&rh���SBH�����"�03I 4�g��Z�E��3�y򞲸�/UՄ��(��"��'�Z�5�[`���~��y���[�ߤC��A+����6Vxl^�4d�cl��Q⯬��d���j��(®�2@>v����,�
w]4�'�8��p��H�����~633FG卖���	��ȴ#u܋'�O�;��kd�$Y�k���1��wQD˭��m�YH�x.�ŘB���6t��G�n��P9�2Z��h<�$=�)sF�!��R�<��'�Z�(��|E5�c�=����]o a��;d�9`��}���,s�$gO_~7����G�m�ߧ�1��q��q`2n����P譖��[uY3Z�.�7|ˢ�Y3�J��e�&�M��}��';��R'=<1:��h�&�AV|�+�C���1�M���a݃��	��}�sg����
�c �-����N��OOg��ɶ��R]����0�A�|���=Z��^��7�=�O �DY�j���S���*���y^��N�A�k����Q���y��WY���ъ2,Dj*��7]�\�9��?�d��0�}dl���,i�	�%=��~�uw����7
�%��>Y
Cŏ����{DJ�� �0k;{L��:���:4��{�M��	S�E\z�6F��,j�PZ.�̠� F��
�8���H֊�1����x?fPX_C��(O�zG	ՓJ`u�ml;�o�A��r�,7_N�c������<eP��1R�C;�8�w[͡���C'u��|_~����`��SC��9��a�e�ϧN�߮ʛ�]���?��T�/�%��J�܆��3p��%8q̘���e�ٿzZ�HG�gj�A���O�J#�)����Ƙ(iy��������|�63 ��e�q��B)�1T0)3�RSEY&�|��G�{��lj�T�B_�U� s���U����w�砜����6�84$tM����0������C������A�!���b������mH^�ً~�]�v�;S��~�'�� ��U>ݶO{��u���㓄v,�-@�}�c��/�o�~3�;P��ԓN
�I�"#�����	a��יe
�E���
�|�4V��I_Ђ�������i�d@&d�8�}T(��LzcwS:u�����Ƨ��������:���|od�4�s��.w	G��v��mOx�7;r�?�3x	�,PXZ^z���u6A�M�[{��+�n�X��[��_(�P7�kvmF��al�� `��<34eq�Ј�<�"f�W�9Ns����7y1���ҥ�js#�����篮��/
��ɇ{��(����b��U�R~��uZ6�������~.��>����$�Z�Z�����P������M�@m{g�td��!f��2�����Ћ(y(L��-��������K0�an��7�O�-Ǎ�rn�)�!�;�u�/1ibp�Ig�G#_I�B�th7���mh���������6��Et|;�'h�=-'��P���찏�lzSn,<4����5�����3�X>�����O�v����[ȅ����m�����QP��yW����*���"�ujO����j���Mcjq)�t(��!�1��+�$�g%qh�V !;�8Cp2�@��Q�F��pr{�0b�ʆ�d (�N�\�s1��'{���ys'�	#G���IP�Q�����e��B_L)��:YI���}�۬ի�,@��B�)Oa��Etro����|n�*m�Tx'5SU���H�'�Z骎B�S�g�6q�����f�/.y%�Oh��mBM1S$�9���Q��ʔ���)�=�f~_S�$(��M�u9���aCլ�Zi>A^Z"P)��/&�0��sPW�(G�r�W�RM�P
��#�F�5+�E6���iCi����fI����ҹ~�cr���G�W����M�*q��x��ht�G�O��51v�Z����` ���<Ǩd˝w�坏�^luE����޵��ޖ�?���'�J�Ê�x��u8 �~�́��k���-�q	l����Q-J�H� \yKK��P��k�Ye�F�0n���&櫩�$j--�`j�X'��e��z06���iZj���K�W�T�̂����/Z�ᆎ�-��>Q�G��!�Ļ�B֖�/��V-�������AKr}m��s�����y@!��������1O-o���G��3�B�!R$�	A�]9�Kk��yK:�C_�)��H�9�8Y\_�%�|�O��:���O�*{v4M��Bu���(�*�>a����~u1v��ͪ�r��`��A��R�w�P�Kg�������������l���v.�@��V�Y���0��=B��M��w�ƺ;#�Staa�y���M@/��0l��*�Rq��w��kz.�Z�& qw�G�΀}j�a�R�it7+������0X�o��k�g�\E�\�FSεQ{ܰriZ�y�k}�Y��KX�?���T�g,Ӈ�mQu!bko}9��#����p�Wը�c�����ڻ���!���`�5��ق.�v�{P(혉�+����%M�M���nn���`�2ر�0�g��P��q�@��Hz��Y��(�5��\�+�-�☨�?W�/���G�.s�0Z��p�_>�q
R�?����-���Ћ�у;0���ㅹǺ|U�N��A'=i�����c��4DT�c#hn�����5�ш�u���Q;�op�uFtou e:��&��ycsK�~)y8
x�-D����#Ĝ��@�����r����$Д@���GM��(5C����(�E�6�'�
g�ԦW{���m��9���ǋ8'�A9	�^����cL��#7ů�_"^�����J�|�u��-f�X-�^���HBL<)һ��dp�+s��mZ����sg��h��.g�A��_%�	���Z���7�,ݨB��3?����wؘ�yW[*\Qu��W>�6)�?O��1��c+�ӳ�M�eN��pAJ�;Yfvf�jk�\0u5G�6+AϽSVL ������@��k�,+��8/|��cY#f?����9iW��^�a���ȳZ�9-P�J�2�ēy2��
V���+ɼ���!�-�t�y1� �����)�&�@gD^��}�a��:����R��6�� y �Sgs��o��Ն�i���)��{�Pֵ����ϓ;�zǎRg�fqYG��C^�����$k����=��0��9:�Z�T�*�-��g�B�	��Y�//;^�r�o���g2{���xq�ܚ����KC#cފ������E�H�5b%?�Ƭ�X����ƭ��{��\��]w\W�/��������޴`\�<ڡ�"N��Y�x��F��
��p���f2����'y`w��5M�0�vθ������׸D�?��g� lO���"�~�E�I���a��懺����~��Qnd��g3�G�n��p�c<<��7��@�T�x���������62�PӴm�]��6E#�����g�r���ǐ���m�(�Z`U�D���rZI��I(���֐@��!��˩]
�pm�
�^����k-�5��Ǧ4�l�Z�N���gt:j�ƹ����{sF�s0��~h	3M�v��5�Q�4��s�ZN���D�9ݍ���ʠ�ߓ;U�Ov{fr��ś�x� ~���u�����KN�mL��O}�՚w�5�l�U/M<���wU���뾻��4A��Lt�q���5�0p�+KW��&[�4��!Ǳ��4G����t��
X�W,�G=�s*Kf]V���m��D]�Jz;�f��L����+[����b���ˁ_����U��ʜ�Np�Ӈn�I �v���^��x�n�i�I>�{r on��ȼ���y�������5�B�䴠��a!�2��eR�^�w�f�|7��q{&sxG[�KK|��4�Y��P�ݛT�=��~^zZ��޻�"������Y9�z,_TY�2.���&�a)=i`D��H[(����f>�9��_�˷���J��i���D�̈́����a�V|p�9ڊ�e0��.g�r�N�T��F�!�Tѡ"\uD�Ɇ�[F`���ٗ�.�(�$&	���~r?��^��)��l��M�(ɇ��}b/Zf�[;�5��bN��_�r����0Zc�('�6�e����wEk�#�x�)��tl�k���բ��������";�݀z%�e����H�8��RN�k�%��%b=/�N��||=9 c���8~Z���B�%Sg�ꔮ�l��H<��L�1g_\��h�����O+�@֬<ٶ�%e\���5S,��%�VJW~�ov�4�=��vu�W�\�J��T��Z��dܳ��_)j�1O��7��b,��!���K�"2�?c|�b!�,!��p�]��^W�,���d'�[����6|�,U����"��0��
�7&c�g�� d��R�-�-���~<�ћ��� 
 $�ŰH�]L�Y��q5�i�At	V
�B�����+O��n�|���V|7-��	�"� �R���Z��`� "+.:T�1�B/z�2vu��^RV�1+@^Z�U?�ȧF/�5��y��g�n�����zhnD��@� ��Y�}�Dxf�"$L·�w��Ng�{�7����֣%�B�y,i%��V�#��Z��	����-d�.�&ق�C�.p@h��}݀��nt��h�����8��X�/<�/�8��������aqNd��4xn�����)��*OS��W�z��;F��k򹰒g#o�����Q��(5�\���F[����n�c�t�Fim��qI�̋Z��P@K�z}*E�>�N��tV9�����L��87��������� {Hݟ��#RdǇ�����W��ș��{uݑfj�2�U��D\�W38s�^��KNb �8P��r�DզY����)BN} �c�T�x9��&gסZ�np�{R�q��6%�U���U�K:��DZ��=$-F�t��}�aO��8-N��>B�� �{&�6=ID�;��.�I�P�؂���]Mf,זE<�C�I��
�D���!�|^_�>"\�j-GM�!�})���<��G�^�NfIڎ����
1�[o��	C́�%�
�Fԑ�#��ۼ�?{��v;��x�G�r{�����Ӕ����6��U�&a7�����������+Q�w�.2�L��#?��$%+eUeR� ��ۙ����;Yy`�$B���`p�ɥ��/��˩��b�a�^��ݰk���������L3�]�Q�5�W�� ځ��6Pm�e՚+]�����#	�򣂲&O��F<7(��9Q5�	�y��428ܷ�A�2h*\�H"1��yf"��{���
$(���?oa��'�B�-J���L
�cުg� B_[�S����,�4u�������3xq�탮>�D�`[��@�X�+d�.e*��稺�ga�p⹪g+�-p�cB?��G��� H8~���mءF	��X�%c܂O��H��B4�0w�3c��?�evHD5����ó�Y��0V<J�ρ�\_�,�n.p&�qķ��BC�9u��w+m�gN/g����P�A��!ɸ�V�� ��6�P�ڄ�X�29h��#c���d��+6��Zh�S	t�(�=��[��Ё�.$$��C��NT�V4��ۿ9��L0	9����:t3'�N�+�f�eޫ|$��#��ſ�G��O�5N�N�� 8����u93�y�ĒZ�JO�&#�{���x]�i�7P��Í������R�#z�}�s��'��2&!_�}�|�PEʁ��r�q���<H��ʇ/�`b�~|G�Q )��ۨ�I�������y5M�$a�����X�E]/ P�U������63e�	�*S�W�ʾY�fS���N�[<Sȟ����-5;���,Q;�њg���~�S[�jC���"�����F{����ƕ�~��V�P����d��ؚO4�9�����	�\J�B"L<�$�E������*��I�J'xI��ѝ*��ō��[~x�����q�C��H�i��8�L�\��{qj����E���(�H�Y7�H U8��I�jR}�@��m�Y�ҋ6�|�s8W�L�h��̉h� F�5f8���� Z�yQ����V?��W:
��琺�c�-6�m����G��{VU`�9���O���)�.��e����6d鹄5�>�wC���0-N��F2��a�m~��;��4$���e��>/����8��o|�I�W�����!��4%���f�rk�ܚɸ�e���}�+����������T�S�/��--��P��8�k�����]F�w��P�0���v~Pvg"ע�E�c%�@hf���)����1��@<��i�9	D�)��we��Bi��`�k}�|e�)wx�� 	�Q�إ�(F���2ވ=�E�md�ݼE%�f���O�G�QH]'8�E�]� ���L0�ж���3#��3�B:ݫ�XC	;`���qy��Wm�d�L�Gg�o�J�q�������8�/Ⱅ�!�� �����>s9�"�NRF9�6Z��VJr�D�ǳ��2}TT&c$��u�4�JD�� ~�O��M��
�aO
,� ZZ^WF�� ���인<��$χע�,��>չ�g��p�V-Nꦝ ���|ж�	mգp3	P.FK֢Crw9�58:c�칒�u+R�6\ԇѧS����"�OvI�6��!�)�\�Z�m�/�@ˍh�i�"���裯�BB�[b�Q���@�@��8C3���^-
�I���B��6��Ю�m����mC/)���=��B�]|_�0��lܜ��Q��khT=�ڠ�gJĕ�E��[�r����i�n�	hq�	�2�>&rM�-Rf��;�}�3����V��U��@&��֘�0��<��4_N�P��:�x,g�q����.�,��!�y�|�:�8����`�d�a���DJ��-A�ˢS���f�@j��@������r�q�{�|����jz�ae�a�p��[	�UK��e00��·�2�yK���;h� Ѹ��F�9��sڔ�M'CU�ݒ���ǁ7��7���M�s�`��[�Tz�"i �n.b����w}#�- ��*sӠ{<a�:l����H�6���RG2�C R�J��R���.Dvl�Z>�����"镅k��D?ڇ
��u���:�i���'+8c�`���k��,ۥ��j����i1yG���Υ�>S����]�h�Ȏ��!��V�����3���z�`��^�G�%8�>�����zT;��� [�l8o�� =ȵw�嶹����@#���F��-���p�AJ���
��"�E�f��8P\�8w& �a)k�[D������mN'2���?�|�L�m�Yph�������
&PW�~B�/+9������eU����yx��^����k����^��3����
���܏:[��/_5/�r��$tI�͚��uF��`y��|��og��C�mL���e�aEs�!g5���񻷌ΐ1�I.�O�t]��0�h�4��J��rH��s�q�,k�{:B�7.��5��~�QG�����OU=��|+�:�.��U�LBJ�O,<�_�
ֹ��t���c}�1�m���Yfi�`}Ҿ6�����U��Ч�&�]\��D�HE�`��G1�r��:uʼ8�p�58_'�! R�@i�[g��?z}�^�*"ah���d��E�4`��S͵�m����8Qn����&��q=�Es馋� �b�<��"�_��-ö�("�3+����)_�1X���E/����j>O����t9ˊ��z�,�=Ї��I'�#�����Dr��Y1���4Vbo�X�9���o#��>ot<��Ʉ�lt��*���x�s�u��j���w�v�Y�:�@�W�9������XiF�Jߛ!�>S���˱���t']�vQ+<�X����F� ���hZ@���
�pi�Y����߫�n�Q*4���S@�\� �@������/��5��ϒ��-P��J�G��{�!�Ѵ?=>�#�������_���"�����1#�K�r]Vd�~�|2�F�9ى%ύ�L�Y�,9�o�A�)��c;q�I�e-,2f�[P`�+Nwn��7c3+ A��t���� ���1��N���Wڃ���<���C���Ƭ���R����_i1x�y�D�{�ENzf��&����9��`���* �)��_a�bp9Z�/��M�D�,ݭ��F|r3�C_Рg�����!�)���W~��� �M�Vw����R
`wX�ӵ��vPCڬ4��쁄	&j4��1���s��W�U�nC�J�Iਅ�,��h��Nbq�D�����\z�V3�P��]�`@�zb�����@����媗��ŕ��>�@%�dʛ#�B���"����	�%1�J2#��GL���Q�\K�HE/���iW�ɳ74x��rc��sT��	ZնO�,0:���ʏTP�^NL�[*�h��(G�2��<]§5�	y���tl�j�`z�o!8�f��Ve6�:7,�E�^�;="����������a��%��}ڌټ^��ih7k{���uO��D�l ��9��m��l]3H=bx����DN�J<,x�W�vZ���;K�G�b������W��
�
�?�����0�]���#o�W�Q�wJq��?��b�D�G�ߧrl��O��1a��i_NL��k�<��*t�����a[:�a@�-��k�w`����7#9�`[�W�Y�K�?��O��Z>4)�?��co~Õ�2��q�N�?Y^qh��k�Z~�rb��g���G/[�� ��nz��z�2+�3}�v$�ZZW��W�wc�*C�x3Z�L�~�L�3҄;�ˁ%��������T�"؍Kr��Z��/�Jԯ"��F���
jL�?X�(ٷ�T��t|ҕ����od�jH[�ZftQH#n��=\�qɂJ��]�L�	�7Zr�˰o7�|<
�h����u�f���/.�z��W
K|(<���x������X��֜�[%��z�aK8���i	��<�a�A@\���v^Q���Zql��u�(�g����ͦ���GW�>� �,�YO�M=^������u3i'Se�]�5��IV�xT���ĨA�*��'Y��(�Y~'rXSΊ�RԌ�����.ZT!6%\���Ռ��@��b�}\�;����5�X�ty����%��_ap�����2L/����=�������� 2������ٝ��c�+	��2Mb�q/[�\Ap��!�H�,p��%ސm2�x[J%܋W�̳�1�!W����1;�Ah���Nd��#Ώ������E����D�{�~�U�@�����{��ߐc�5��Qyׇ����<V���|Q�s���jl/�=̚���m:#��>~;b
3��������r���PiBIpA줣�nT�+|?�` �ǍX `U��T,����jܻ����+��2G"{+]t���ZoNw��3>��
7�ٙ������e��r�6���p��"�=|#�1YR�����\�4�V�)k��Ok}1K�?��+b�� z�YЯT��$Ixe��/AVN�|Pm�����C�DEA#���{��i��,�)H!�6O�ʓH`ĖY�����T�8 ��9c��6q��*=�aʙ6gzm7�Y�	������hp�R2�gak��Q�U�1T�iy�Sƹ��t�|���F1�U�-����uC ���O�Ļ8^�y�΅w�.�W�I��Y�y�F�S^r`/ZM�Bc�)y�ֻ��ۻ��A���|�#�u�^�X�Zu�h � 4��Z�Tƀ��J�c18��k��$����0Ff�'��5�x�p��^�/��.���,u_]���|&K=���=L8�$���wZZqx�4]cp���9�3�x����R5���@��b�t��1�7Y�_&�D*i6���٫w�"�U�I�\��x/��(������a���.����Cs��z�8U���I+��B��yC���j��;�b\C�ٳ��ޒ%��T~�lEc*fcͨ\RI����5$�}ThG]�0���z�BmS����:�P��eQC�;�F�E�s�2��r�F�Ar��d.V��X%D��CXlxV64EB    fa00    2bd0uB�����M!��g79���c+��@��;��%�'���������J!������M--��Ho��<�kŇ�4���j�ɾ)QZ��<�.5�nQX-t�0ZN�KZ��nQ~AǶ���v������]ٷ��Ԡ��6���s�/f�a���*������oI�U�ѡ���;��p���R�I��(�|]7i����lvU���;=/��pJw�O2���%^즶�U=p�����}p*N�5�\��./wE,Κ�!����\�f\��:�)��L��\@�$��-�5GǏ��(��H��3���a�^�����6�.З��CP��������m*.��,A�O�DZs�oC[�������ˈ����fs�L��G6����D<��%k�w_k	pg���v,��LCH_�D�%=�؆�k��
�er��RK�Elar
�vD5�VS9��	����0Z
�G��ޢ�9�/�4N�[����A��O�֢ɽj�;|".T�"Tݾcc3CԲ�8x�vI;M5���ʿ��n;��+�5�Q��?rB���M��a�u#���7��#T�!|�`j�~��s�[Z�=eK��~�L#�#��8������><D��ϰ�:���� �P��4A]�"����T�6����9*�t��*r�~%�g|�}�%�����)��d�-�S=�Y��cN���b`�S�'Q���������z�.A;r�X_�;��PX}b�����v�=ki����x�	 )"+@ņ�:!��#S�Ý��w��u�����E�w�i~�����Y�Ny;L�·| �Z6��I,3��f���fV�3�o��X�J��Dԫ
X��	�����~2aB7[i�(����l�[䝹���;��Q�tOn�\,y8̷��\c �fS?�@Ч��JGY�5*��И��{���Cl1MM�C;����ymyh��G�-G��A�i<�A��x��4V^c����:)�u�>��`��o�=O~�m,Y���Nҹ�l�2`����K�d�T���g玸�.��w(��i�b</���aܻ�R�I>1�9����vI�r��Tϧ>���
m��Ǉ��ۢ���d�MUblNE���Tt|� ]L�a(��-1x|	<6ԩ�	�&-��U��j���G`%Ƹ����\{�`�n��<� �(ɴ�^Wm�����u�&0�r{kU�1�?S��}�E�z
��+|���_�����-<r�al��[Kc��\7dn�F}� �05٪���,��f1<:��5���U�8"ʅb���	_����>L��U�Ϙ��8��k}��F��8��L"TAk�*,g �����!�Țv��	ƶ�>dD'��vp	�koj����Bm�Q��{�A��=ͧǤ �0/�v�S�ȍ��&HY����)��:Ώ�6$����,M D�x�a�ɶɏW�:Rݔ�O���0�9�6b����M$�Zq{�u�q�B+�8kH$����	�F�<�B���]d�S�XR\H���ȧ�6�3�&���x�Q
pvq����S��-3�d�?�����cJ�m#u	����v��E0�:��&�G�[fl���1J��S�F =!U��\��;\���=���%�g5l��.�s���)sp��Y�#�z��=�{=����aҳ���VdQ9G�*r9v@BV�	r�́���!�oJ�E�N��,#W o{�TL�i6`H�iA:Nɹy ��#Nλ[��퓪�[\04��N�y9O2�$J����v���|��t�5�_��}E.�R�0�Mo9��d|{1�7��Y�{S��+��gcg��:{�9(�4��z'Aw�t�";l]�5��!���T�39�"rA�.!e"�^!(_Y	������p��6�/G�����Y�F6�S���j�n +?�Ǒ���h�?�d�%�}���1�nz`ߒ�j^��4,�H��jUzܠƏ(�A�r��FS*;��
嚃n��t��^X�F�b���$�V�;im��*�_b���PT7]<��?{�*���g$��QQ�'��� *�􍡼�1�}@���]�XW��5���J��
�;zc��V�"ы)�7��L�G�8e��pj=�U*����G�C���:�N5�e8щX�g���B»GB���v�S�!I ͞}Ea�N����8��Kj�u�Y�M����x��`d�>>�y �?L�ư����=�;�]+(MZ~��]���u�G�gC����0����K%�-�s�%9��t���r�o��J�k4��x�b���22�3N��DS�6��c�|��- j<�C��2P�Q�&k��le��.:3��3e��&a# 0����	� �,�N\-�^�)��5��{�Dg�.63O3��I�8i�~�Py���?�KK���!_��nt1�Њ4/涋�G�]w��M���=68���T��7��.ǘ��À���Y���t_'���=��Y�U�YS�Ngc=��T��9��VNԠ���@9���c��-~l�B�/C��iw>h��&J#;[��m�~�[שHvu�uäS�B��R��:����e&��.k-h%;H�~�c�>s� օ���\��S/���\J�uV��p�Y&�bT����'lި�{m���ވwr|��غ��F�!&W����ْ��f���_U�ti�[¢�b�"p6���O"�t�|/���<�aaz]+-C�\J�[�����C�Ⱥ�?�ڨ�yTv��$?ݜ�k��|n�<��k��/Kh_�P�C�P��ʿ���e�د���-�������G���|\.nvq�Rq=S����*��b���{�/���OCF����-��Wl� ��" y����?3��[�gY�!R�82K��^�-EW��ƍ-�8X�!�>�rmx�h�F>C�rVi���W2W����ЍcD���g@��u�����Y+:�*��T���:��)ӝkvYE�C�y�_CO�g�����{���/�lm|9�M+�Z����Ǫ���L��+�jU`�[�D�A�|#��cl&L��V���[i?���u�h��|�Q������=�^�z��F��2�6]Id!��WyН��㫶ڍ���?��V�|Ԫ�9C�Ż��U��I����c��w�B&��@�R���2�A�����w���ʉ]ݚy8`
�&�o��e����ZQȎ���mD�TDeR35/ca��lͅPF���$3��@��b���Ӥ��j��1Z`�v����`�V�p���-������ࡓ�̼�ȃ[�i��hwWa�ma��%3!W���|rZ�杙��R��h$�f�T�e��rp��;���%�B_]Rb��#3ļ���9ʥŐ��Ŷ< #-�A��Q^�~��7q�d<x+�A�ER�α�M� �\���fi�W�xv��x�Xr��Z���{3��&>�S���^���b��0��^`r��v��fq�&��Ԉ�OMV��#�4��t�f� hP}��5�Mx/q~8T�di����l2�H��髻��n�*��ycX�h�6����1����K�qEc�m��P��a)x�؞��/��	�;}�g��.b�@��n9�ZLz^���<���7pw���R��vX)��o�z}vva��	}Ř$�o���}�cVC~��?����G�d��o�V��YZX~Ǵ�q�Tk���>)��Jƭ9�ͻ
%��R\�е�*U�I8M^�1;HG�fܜ�۟�u�B��t�<�:�l�_q�)�c(B���U�Af��)��zʘ��0G�5����F�U�A����ЯC-����p�iv~�\��m�m&e?ҼE��ݮk����v��_,z6�K�n�N�9���}g[f"��R����(Ū�ʢ-���S�P���֤����� �����h=^M�Hr:�wE
�ua/k�H�#�4�U��m��@a�Y��I��H{y&�#����,�F�nq�}3��g.�&'?Fq)���'��Um� ?�ap{�.�Aۋ��:��\2�::�?^ NxOcIEڌĿ�vQ�����/�)J�c�b�)�m��m�ዡ�ը0Ϗ|��W��Xrϐ�	_���WZ�Ҟ�M+�,:q��}��#�����	*p�(x��_�c������`K�1�����q0��z4hv�6m5cԥ����G��$�S)���|0�
�o���r����5D�ENu�݉���I��� ן>�;F��ȷT���[��h׻%�R_`�/��2�$��}L��hMX�aNO�A���#bN��
!��O��9�i�3��rQ�>�鉈�MJ15#��
Y_��C�c\��I<B:d,;�x�ƯI9��,5J�3�A�؟%�kw4�4���oY��k�C˭����X܄�5�tsZ����E��0���5�e�.�-��7湺1�= t���ٴ�Qa�T��W�s���AT/�>hF	����9�� J2>�b��9F�Y������)��d��z��wJɍ�fk�����~���cU��~��H��0�h���vFަ	�o[�Ѭp�9�;�
�pI�'P����Ȓd�kB�����ڤ���J�ծ��0����!�_�Z�*Y���_"2�����"`�3�j,}�18��`PL�����]�)�ӄ���ڏӢM�D�X�ttZS_RQ����}E��d�d	Z�<���a���a����F�O��H��)c/l�Ac��f����K&s����0)F{�F��B�:euuFZe�$:�� ��s̛M�\Bc+\�J��쥳Z�a^t���ܪJm���_zs�����"G�c�g�w��
F��
�F;!c�@I�x����S��(�D8�%�cB�Wy J�C��)�6u���9}Q�V o����QK�y]я��q���;C�C&�4��Y�vr�LKeŏ�д��
�Xn����.�p	A�����D�m�. �qS�	>��;�A��߁4@�#�[�jjN�����ê��eev����y�s�~��nz,7]U���Q��@���V+��W�
 ��#��O@�I�v����I���� ���JB$ܸ��#&��_��eM�-`V��v
�=0��A����Z��r�5�^I��ճ��^scEz�W��',�UzҒ@S��,�X��O&
; ���� SC���ݸ`��dIS]W��e}�s��MU��L\l��wϐH���(>~��� �b�%kk�n�`�*�2,h؝��7Wx ���a��e���C%4�!�p��k�O���q(�E��&�o���@�ٻ���&�U���+��&���1tW�C
t�<#=n�XIr�� 9��-�ȫ��%����P��qF��T}�Q�h�֗m�o�>4��V�?�$m��`�g�ﴈ�i�"Վ7UO>ĻUϞZ�䉆r���m�V c�L�h�'وd�y#�
=je1r1�A���<Κ��:��@D�VM������{u����m��|���)��s�|ܫJ�I��~FsE���'��C���⾃ ���
�^鄒���$ %�Ǉ/#5?��QIF��p��޼_�h��"1�	�H]uL��~p~��黂8!59e_�@}�L���|�Ϫ��v
����ݰޖ��}%���k	���W��uS�@=[ߎ ��7��"=^~daS�k�D7b�Xtxu͵8�|�
맼��̌���^@K�X��쒿��R���G(]\ގnH{�vqﴁ�ϧ�[4��X�O��r� ��ߎF�t�|�(e���R2)4!}���tS	NBC�!%�ݦa�o�1�����%�_��E�i�6�� |� ��8�ea�(��mwX��G����g��Z���hàu�jP���xJC������ �$�q&}���'�9Gq���c�Z}�E]���:u�]���ȳw����a�vw������Y�l� J�Lx�����	��W�BA�}��SvxݖfA�,;�qGϞ�x����������ɦ��o�_��=m5�6�#8���+Z�_z���\�en�}	@+�ڞ������)޺���+�I~�slbOy�3��6�zO=N3{���_t"�؏�nv.����SSF�Pb#��2�������]��\�� ��g*D�ZE@(i�X�84�W�4
#��")Zمh� �������d	֓�A+`F�LOr��{B����Y���'��-#P�1�V��	g^��VI�x��=�#�(�]W�p�݅�~��G�w�?�+t4��I2k���r���Kω�� D@�hF���4�*G�Ê3z@q(ם0��Ų(G?屷0��[�/Ҋ(ɍ[�|��d��PB�%؇iRe�"7|2���´�/��w��:�A+��:p�M=�v*���W��g0]N���̟M.JF[�d8�{��ry�N���Q�%(�as��
^�
�n�n�#A�(3ǊH�ݓ}��A�#����ѡ�9}O���Hs�8�G��1��Gj�t�Ґ��U��g����T1
Ǟ��oZ�MA��.�.F�"$�����c������n���U������ /���
�]��V�;�v#c9(J��ے���y&� �A*�k�	V�1����@��Y��y�M�(#�T�7�y��!��p�s��lx/����)��ӓK6h{!�/y!��a�x��
�:�A�\��O/H��8�A��8�&�E�5������Zv)DO�j�pz� �s�c���dR⛖_����Ϩ�����j_6��k��x�\�zD
����U�<͎be�7rq�K��̪������ݖ�!��7����l�mRCSmyS��G�\�b�f_�'ƿAkzn���~�Z����;A�B7�"���W�'�͘yVy��H��ׂ@�[�2?%��_�\p'Z7���J��Tf�����*�%:�\�������f�5Q��z��hћ)u4�|E��� �H��\P(}��4r�ϔ�9���ceRYX���1c�#"(��x�џ)p�x��Fvy�f�O3 >�2��F��Cxs��aYD���ߓ,�M]�4�����o��Qb�0	C�$q�P�3��L�#�5E��in�<���/?Xg������G���d'��u����յ�W����K܄�Ç���_K�ܫNI��ɢ+�����΄A�(�T%\�����%�B���Φ���_�s_��q\J%ܲl*{Z�\�,r�a7���4�f|[IC��n�W7�k�|��a�>q�o����Ǌ1��1�b�H7I�j�[�HV��������%[Qn�`��!,�2������B��
^Z#���#)F�5Cf�jQ�I��f����P
������w��҉y趇 �*�Ϟhժ��7(s(�1�#�r�� IP~�V�xV�Wyk]�����f���F�$�D ����H���Rh���v{)��m�/�oҍW!��À��=�����(3%���,�B���CR�=��x�E�~������w��Pg60�x�do�4釕=�
� �kG,�oq�1<-�X���m�q��e�����Hǜn<Ζ4�*/+oЈ2X�����_)�1`��?ew�*ȜU� #��=/1��"f1��{��f.'w�A���c�X$a5`7�B�:�D"�4=�?<Y���В�S&���a�Cp�-���s�B�'��|l�
퓼�Q��!b�?���1�`�����&cO��Jt�1bT�V�_A��ߑj5�˥����אg;�Gό$1�A��Ru�Q������x)�߿��u��w��,eJp�z>/�K��"�6�X�t5b�vykO:��謚��\�d�������&�@G���/�͐$��/@���N�{G���M�6��3
,�3��s̵ X��wI��B����+ζ��e?A���� %��x��h�L3w+8�M�MS�/v;�A_�6m.5�5h�bkX`����q�M�L�Y����>M��|��v��f+��tǀ�|�H�z�~�1ᢠT��j;�\n�}�Z�Q�M�FM3��e ����ѯJ�`a�}<���%�*n>�]8��3%��	 q��	7�lAR5չ���zO����k��D^��Ĥ�����">������2��lX�R��*�G��? 0����D;my3ı��J$<3M�V��^���D�Ҁ鹧���5��X��NR�H �v��o�Y����Ŭ]��Q8������$ٌب͍:�-�Z�E*��$�d�ғ�-&�����	Ө����T���E�*���/�; ͓��:<A?)�Lŏ^Ą�m}���"����9!� '�2 C5�r�|-����gIHD�<q���S�x$�RE"�[U�XV���P�s��@A��Q��M[7ئ�툣i�%��zc��e֠H{E
[ۡvNQ��
�vk3����v�ahV&�e�K�� �+�7׆�O?:�!Ԩk�5�kq�kı���q�or��
�#�$���M�p�@��EvF�)��������Z�g�32"(����dY�d�?���x=j
�*B��+v �NG����j�'J;��t2�c��y���b�|�VErB��J�,
��w{a�Ք�n�b�g)����N��*)�ܠ�ĳ�Ր�6=�>��w�� |N�-��)��BJ��y$�
Ѳ��J�u)����Z|�=��/�N�j�Ӭ�Z�to��%�3]V�IЏ��_ZA�B)\d��W	��Wp
�p����P�+k���4{��a��4Z c��bvH����xU�L�MS�;˨R+�Ĵ�����J��e��nҭ-'�D�ev��Y�s&63<�,`���L�˲�U(,�I*�@��\�S[+` �����	���o(�Zt���#˄ěc�`������>id��ظ�� &�#*ה�D�v���E6H���r�^�1Џ�u�M�!\t���I��}ņ���כa ;1 �}�
��W����D�ⶾ&Qٵ��.5䂟�M?�޵�x{;Z��K�+�f��M-��ȿ����2����� �A��`��N�m[M���!���}4��P��t���4�K��'�+�tzה��?]�<48�kV!A�3J���c!��-��˖�%"
�xJ���/�
gꢱN��A��RPx�X�VЗ?� D&����S՚�?/+Ē1���d���Qbra�'�i���OU㇋h���f�3av$�n.���~�S7w:�L<���s]~߃�7u]r���p����8"'r]��	��͞�6�ۛ���(�-�Sf�|�i���b�]�⠰�����YsZ�:%9�1�G����Y�a5��:� N�#*N��n=��K�g��S�ES�P�V5���_ezNӔ�o��[S���<���e�Q�Ҥt��IF��C��ܽ{�3o`��r?.�X�(%jz3n	�0�O�ÿr
�V�5�}6p�ڣZ<-ǐŃ�JKv."�=v�7��S	�:E���j>��	%u�vf��Ir�Kֽ�)��}�3>sj��Q�H��B��qq-kB�\������s�ыw$��>e����G�h��\�p;k�U~z�4v���aVØ���Vv�J9\���Ƭ�!����">���!R�y�C��ߠ1(R��b�ItAy�rO-A+�eCB�z9~�[Ć�c��f3*�L��"�����ׅ.F�s!*�lj���Aݛ���纈d��^%G�ܨJ^���4�(�����/Z#�2�[�`7�NG���-��Ҹ���ۋ8	����g��W�v�
��%�Z�u�1E7j���m ����O��P��\��V��_�L�MoL�`����9@\�s��.�%��PjAj[
V{}�"R$���O;`��7�w�%���1���o�f�븠!� ��k�P��g;�M ��f6�K�?s�G���iwz�?k���3"1BY{%�0'����z,��~?�헩��t7!	��Fʡdl�7n�J���n����e%){'�Z=��b|�FY�9ˏU4R�^vLZd_�܁��C�_� y�S�a.�K��ϪJ�I�V�8���x�����琾��?���d� �(�Qq�^~��D1���\�͏�c�m�Gß/�I� �J\뒺�$��ܗ&� ��U�#�,wJ]�C�#��S�161yN�z�К�K�o´�@gx�2�D̸��z3��v�Z[�쇓�w���p>Y�gG%����L�?�zH�k�ÿ|���x?2"��`�穰�Ao�:�~κ/V�T[�p�|����-MC���؈Wɳ�l��AH9�RQ�6�0�n~�`��i�`;8W��\�p���w�ʨ����	ۍ��)�_'Rѵo!�[�����|o���ƏD!�r�����>�Ғ~�" >	՚'{�N��Px�"�"8&Z�>�7}��)a2D^�u���7!@��˦�C[���j�&ʔ�\κ %���&$�[����W�'���`Qwq�,<��z�˸(�)��Yr���cG�k�.�|P�g�K�Ɉ����C��q+�Ux����N�Zá�^[�c���������D�:;�z�?��n>��)8wM�����u�t�?���F��Ӛ����^X�T�)�/�􌈡���y_��^���g��fG�{+~'D�Lr�vw����k[����B�u���������=s�_^�Unn@Ot���f�m��;{!�&�9�jE��5k�K��[�Zk�3>i:J�l�B�����FÞ��<���ei4�X�F�E/۵�r�D��i��̌��e�.l��h�Uj8HJ��9j����k��4^J
P�o��,�1��(��a����en,E����з#�VӨ{�JW�A��y��-@�'����/4�؄�*M����wwN�<�{�Z�?_�΁9*l�mF��X^�h`�7R���c��])���_iݴ\^�]�!F�\��{`k����)f��$U7jq�$�ܧ���n���ܹ����%��;I:z������(Bw�����ߐN���G��Ǚ��Z��إ%.�i���|��$�B�����v��R	DFSj�Q�G��R��%;$Z�`�p���C�Wd��1 %lļ3���|Oqj�ڹ����!�Xj,4H��>Tk�A{��*V���e�}B�;����0F�ԙ�[x�[��ԽJ�����<��XlxV64EB    c829    20e0�)R{q�S�|��FxhOF�h��������{�Ɩ�~�nc8���7�*�a͕��5,(aє�L�Zó��╬Kv�\�:´����`[\�Z �F���T��1�k����K�~0w��q4��JF�1�FT(�3G�(5���"l-�=�\ϣ�>�XV��5R���Z��s�����/N��{-�d"+�@��!�6���TÅ��~�;Ё6hI?��u�*�O2�<!���ۅ;���=	�fWڷ�i�	�m�_�0��B`���n�{^����i�%�>�='âЪn�
��3Q���T�ڄ��&��9vg(�I#j��.�}k}^0��]&7˓��&�f�rE%
�&����7��ۭ�A�����z�~+��k���56���:��!�wO���(,��t�<Q�KoY9S���r������S����JP���eA�GL	��g��9�O�"�'J)zе�F�yt`�����rS��?���L�.�~]̔�n7 O/�}��l�_�$��ۙ��ȷ��W�5�$v~����Q.dk�A%ŝ'��ds���):������/�Y�zwg��4��oޭ�ɜ�G�}��F�by�������!B��OsQ>�L�[ �j�GK�v�m�Vt���.
��i���=H���_��3��2�����1!�a}��&���Z)�=�PF�����CK��ccʣlm�0�S[����87(yy��i�.�O(�$Y<췵�иAz��o����Sю�ō&G�ĒX�>��Qqŝ(������{+����9m�ˋ�y\K�p�pa�z�Gq�e��i.#|�ض̰3n��K����%�.��[�qM	�ݚ}?z��}��������6�	��eg��O���x��B1(SRo(�`��A�6%�Ǆ����o;>���6$�J�9X�)�	рY�[�B��"Mqo��=���k�-/ʹ�;�*	���P�(��LH{���H�f�^���@���čN6A�:(B�؃ �eqE���_�d9��K�*�x�����%"����1�BT�_�$Fu�l��9C��۵��~��XI$^�ӽD�)���69H�s췰3�]�kG."+?6�P@�Cd���E�^L	�EКe��|���Fm\�ӿ��d�3eH=�9/Y����xg~�L�$i�U��9w�>��7x����7�VM��n�~�I�mM4{�Ukp���"=���/�9�ETK�l�߿C]�l }�߬�^L,A-vʐN����j8�LE�W�
���n��ă߆��������>����liG��t$��'�'��#Ȩ0��C���it��ܙC�����d��}6!�o"hM.
=s���B̥�w�n��KӔ�O����*�_���$���y����`Xߓ���'�w9�w_�Æ��;nI��:_:�.~���X>�9�n�s�z�-����Ʋ����ٙ�]����}Ln�^�vM��^���l�ռXTC/�e��Un�����Jat��ց��f��F�E]��k����}��ШY"�-H6�ႀI�_e	��3���b�"oK�6�=�A7+6�V�8���l�y[��*�ʀ#�alͳ��+��Ӭ�:���xT?����6D�6���K�N��]��p<rn�js�����5.��6B2�87{�K��}2�b ���5�)�����!���{�ʕe�""�@kҌr�	�]iiiK4�j{~���s���@�,��p�}w!S���n3�3�_���&T�ل:-��(J�����-T]��x.�l��T��;��3�Z��D}��$OL�	\q������`;$���쫺H�>In}7n{�2+/�W��9^Y�}SޜY����\Ӷ���d�{��Ei���������%� }��Z��ޡZ(]B�Kn�\�����Ue�A���&=�Ҹ� ���	�	���u�19K��������t:q{��^�m�^�\h­�>�G7�CH���VZ���C����u�{����7g�I�����h]��j.%7�$AFpc| �ف��Mo��=H�.Dŏ��-.�Fn}uy��^n�B^�խ���p�Q��rHt{�~�O�4�lc&xG�g?䚧��TeB�LZƮ��$n�@-v������>k|7�`͗��C#�/��*��n㿘A�\��;\W�E����%�FH��LV|�E�{�2��~�)�`x�t�t���g�/ޗ
|hk5�C�#�(��8���}$���V�q�LV�)�N�X�����|Z�ӏ�
Z��49b�W�(��?c�� �����!a*�.���;h{\`S�.����6�`ͭ�4$2]O�\����"%a�(���$�3p�櫍�C�6���h�N/�b����ϕI��Ow]�(��Y5�4<����{�?{e��(k`>>�x�y�������ɧZ��1���1�&�c~���i��9|
ң��&?N�6�{DW���}�28=+JWk��#�I�>�;��Ⱥst���"K �2v�#���7Bep@��F�|>�P�P�܉`�{���~�p�C�Sd�D�A��G�,`��~��o�]q82f�
�(��ʥ�?!:)��U��oռ3��iI�[�OЪ��a�ދ]{B�
"1 J�)�!L�n=�<`MY�o_�����J�|
z��)��Jz(�����^��XU^�-���0��J����ZʃՌ\-z�muЍ�yM�?�����t!
 A?���ަ�wx���W��Bg�N�➏w�A18�Cg�6
{� ݩ������5k�B�v�)�AC)o��|���U��U)#���j�>m%�gSUx7]6��'A#g��R�(�g0H���Y�,�[���\�CĽ	!��g��vry�W�{�h����3�?f6��y�
��7�9]s�<uOѲ��J���[������*�z�1�P�W��Z�?�i.�R�8��;��@|S2�D����X[{�_V�ơ�K#)�`��4DDŌI�X沛�{�Z3��	T�pa�)���v����ɳu�!����a�ֲ8_M����"(@J�������5��$�,3�l��>�{�vu�3�o"�w/ȑ����a+��.`��
7���-�\����9��ҍ ��+<9&�=��MJ���|�}����9!�\����h��S��P^�w:�5, ���A��x��{���:7�5p��%cD��1�?��z��/�k��~B�E��Mooem�&����&#C�s_Թ_�'���	��nY��b��g��E����ģ%/�k���ܦ�:��{93<���^bhd���~�,�Q�����N��jZ2O�i`��xN�9�w��~���w��|%M�S�E������.��
�,�j`�z0U�>�$=
��<+��ͫp�{x�>#q1�����*Qm].��ԔQV�I�_�<���7�=�P���
��oy�����GNM
��P����3�4�6%��Gr��o��ôH; zЛ9[}\Xe��$��P2�4�CP�A�Mf�}�TW����s[���v1;lj~-"�i�S��b� :�Y!���~��8�_C��_ �������ۧ��?����ѕ�C�[
3���f����F0$�G$�m��u�F?���{�p��Wp��H�[N����0�mc!�!
#{\汭/��k1?�����1�Wh}p!V( ���2˦�JQ7*{C	}E���ܣvЏ4��i7�;z��h��^�F�W}���
�ub3$3��~\��aMÑF�͊�A6mG;�F�ol�\������r����N���|ZdqP�~7�}G�v��'۪������B���f&�~\mtYo6(���1�S������.�z�p�؛$�c3x���7S|b���ó��~���p�G�-���CL{�����m=w� ��4��������=�q�	5��X��+u�D�ܦ4t��`��(_1N>�x崇(w"�^����NX����Mj�u��|�C�ce�{���6��H1�П�s.*��p�k���-��b8��4?�i�z@ro�����;@+Q���dq��B�X���������hq<�8AǪ﬩k�][K�0�St�\��v�Ve��	��=�QJ��w�ӿo�� I���C1i��d��j�U >@C��+N'ν(���.�vP���%��U�-�A�@�������c<_N��}&il�j��4�X�W��l�]�9�2����y|�HG�^��#]�)j�'&�퉸�~�M���h������5�������L���F�T�����w�g�#�؋�E��C{�� �=@����v��1_������`�=�NO`�t�;�dC&�`�B#������L�^kJ����'*�7�
�"nJ�4k��k�-��a
��r1�r�*fPA�A�"���!#���
���p���e�!�i?�ܴ>3�qt7�2��p�Qx(]��Q��i�A�w>6�ĩR��C�4��2��L��y���֪#�Ӣ�G��J[ʡ,�]�k���L1��oA��?�5TlL�un �����O��3M�d^���%�q�6��){&"~���~���Ѧxɻ��2��d�;������=����q{x��Pw
��6���IGAA�/~Q��i�������/{@��v[$�2�J�U����W�/A�'l�ˮ�AqJ��u����6Z��ޥ�Yh���$����Ԕq5ts1.qq����ƌj$��F]�2�;�O�7ߣ>����%EW��@��a���2%Ƥ^2Y95������O�/���F[���&�#�C�%~r�d
N��=R�IK�ߞnf����=5��j����b>p��5���dF��4�U�Ǹxk��4�3��Hɻyh�X;�~�&��A\'	Ɇò9R�"�&�I�3��i7x4�c\癀��#�Q����7�j��=���،>ޟِ�mv��4��d�����{n�=y(Ax(D��ѥ���k���❬���x�}���}�r�임(ތ��ȹ�ƙ|��en�@9Ywz�U2��v&��ax#��p����)��d��;���.��UpOѪn_��q�y�ś"��84h�-��*�w�(p���}�&���A�J_'���Ck�#�Fe����dTV�#µHî2�Ƕ��K{��$ϭ�8�GW�g�ն0<�l��w)��u��N�&f,s6��p�a�G6btw#�U4�2�r�GE �CN�-]nܹك!.�QqA��6�~o�6dy�p�.a�o��^�������+�ƘF�?I/v���IV�P����(��"g���e�R��� �^=6�~�33fq�V��^�h�7�ŶVB�%/)��)WM���c�+��ev|�c���ς����kX5 ����52��ꘙK�i�J��/=n�*��S�k���o�}�5n���?�ah��@.��R/�.�/i� ihG-��Ŏ�v?b�r7鰆!��t��W/�D!Z���+e�K��QDl	��ߩW�
)5D+ctP2��&҉�R0Y��bb�Г��}>դ5���9��b��,������0����-�$+�@y�>��&���\k��ߋ���c.��ۑ?1 q"j*�"���[+,�E/foO��ԇ��6IL8�E[:!\��=���v� �
�J�]�ؔS��r2*��ȤI�/��^�#��3Hz���(q
�2$��>�rtn��qߏ�&+�M/0YN���r���Ar���`��{Ŭ��-t�c%$
G�:Z�f�V��h�'\O>�#[���H'` N̌��{����v ��0Xo,�PJ��3���q��{����O���'�O�=Ke,KH��ɭ��/�;��s��jŝ(M�¢/���.���Vɧv9
�/�k���t�C�AJ�������q�����#���0E# 2b�O��<�]:ӤyUqy��5��|�u`��S�9y4�
���5������2�(�О<v@�
T��%��t��U]�g�Z�G��zy$�}J$���gi�����Nm�ThB�^�������X������	X���P�b�b��b@ׄ�a�-���	&8��t�v'�\`�mX|���n���jmw��pı�5�X��ͮ92�E��@w����c��P�]�C�F6l�+z���Y�6�x�	�����ybJL�,G����~�>��唄jWLf^'HH�2ZpA���y8��Et��p$�7��m�!L&��}S4�-s��p��{��I_tz�R�n7����e�8�(��%:]�E�6������_��΁�o�w�('Р�d��/Q�KQ��d>�L�Wx;9��u
5Y-i��}{��������*@-d!�g;"���x�Y�m#���T��a� �[Nl�j��<��x%�nHG�v?�""'��W8��M8���j�+���4ү]��,��R5�~Ț�k�*�� R���.t��N?����>
V����$�i����A��2=�Fӵ��U�����P���e؂�"h}�%F�8�4V2	��ɢy��5��3yL�Y~��ݬ�r{��@�`�/3ȻV#�ʾ߲n�աR�ɫ �2���C��Lsr���z[W��qE(�Zr���F7z��>Q�Mz�]�����㡩H`�'r<+��.���"o*�׽h��{�&	�7�l{v�~F��k���Uz�Z|0���F��f�ت��w5v �
�Vi<�b�u	n���Cz���R�ȂI7,W��w���U������Q� ��	5A�]X�C�as�5ե�3��֘��X�f�8���;���� �x�Hd֊�H_;�!ƙ�����B���H���ّ�IE�J|�━�}6��R�rO�?�Ws���7�[�-�Q=�(�jfG� �N*������I7e�e\�'�m�h�; ��ws��p�F5e��2t��^׵�-��'�Jl^���0���Yy��]!T�T�V�Va�x#�:H�&C�\�[U�ٞ�F'V0-�f1��]�;��z	�^�"%ch��!(,8��f닀܆��s�v��x����#��o?��3�b�R(������z(df1KbW�� 
�V�K��ln��D8$˧XEs�?�����txH{W_mM`$��͗<)����j뼇t���
/��D��5��ds,kY���o`�)g�T����.-5����g�*,���>>�!��D�j�i���2J����C�d���LD̯�D��TfM` M'���b!�����'T�Մ=�il�屰?(1��L�.S���1U��Ӿ�[!<F@��-����&�R{��'�8'5T�
�h�����%���?DL�c>O�W�#�Y�b���>�B��"6�גC�v1�5K�X�<����J�y����`G����p����D���P+7�9�Vð�p�}�)�&��YE��Sy|����S��]qB�S���%_����MCG1���.$��G�t#7�T�@EQ�9	/�y�E����^U�tb��r@ce4��īщd��������5����*��#�(5Z;&JF�'�i67
h��S�Z5�[�� ����"'R��_&�5G/<-sݤ׽�$��y���=x�oA�/�%����0bO7ʉf J2����z��F�������0c◔�<sBR����5�nz�&�W|.|r��P-RI�<*�.A?׷�L�r�7�2Oz���O�h,����%����3*f�I|�F�V����"��hrY��R@�v�l��.�/� ���/mFx��
��V��;��pM�]M����m�����#���9�%_�B��)[�۝VPZGoG�ɻЗ��L�ή+�}w
��J�w>�qŇ� �s��I��[�?c�o� ���t"�1�pW@nbd0��27�(���
Zܤ��^�J�K7�`�Y�oi��`��SY�t�=��S��H��`i,������*9`\�s4�=�ߵ#��7eq�m�/&�r��<G`m�H�1�y�av)Qn��I��w�u��[7�7bC��G��)�M|�	�l*gN�0�[��Bcנk�\���/�i��QF�-���0}�{\��S�s�����Ta�HMo��pf?�CF!��v	�=�y��̑�vLJ��P�C��|X��/5Ҋ
�$���F f�6(Rǩ�H��wtT���������ȓ�ѺZ䨒��P�5�]9:�5���&�ޜ���F�SL->Y����G؟��n�J��!ą�&4x!-���驹f�24��	