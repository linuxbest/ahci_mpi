XlxV64EB    2134     ac0��k\1����}q!W7	����v��)m�zJ+f��ddQC?rm�7���H���,��5��1@�{Fm���T�iV��a7�=p��JLM�"�T�2	�GXS4�i�|n��ÄS��L֥��Fº��ͯ+��<^���L0*IL_��R�m�$i 8�*����@a�?�
�0u�1�#v�a98��ШCZ9��.R��8j�����������А| 8+�r}�<��XAĚ��\ռ��Ab�\ua�r�3�*�9�.G�@KF�hy+�*X*܉`�&zH��J�x�p��RR�%������'4bj1[;��傇�A�R�w�$"<qd�y���� %k���Iaĩ���Q F�I��u�r�L��K��1i���gn5)�fdW���&�lk.q��	��D2ĵm�ά>�42�V��ҮA)�J�{�M<f̈́Q<f��ִ(ר�����;	���V�dn͡@��n
�և�09�r�7Hr5�ad�릁�dQ\�(s@��Q\+�+C��f#gĞ�dq/���QA^ ��^�JC��3O ����Mϙ����9v�dD�5���*\\�>rZ�8Z���%p׭mogt�϶Dÿ=ę$"Lѕ1������r2�v�T����%��s�0ُ?U��"pz�����V_�0TyT*V�A!�f��e FL��)q�� ٳ	�)�Pk���Ix܁%��[揀�	�qN�0/�}�z�R���S^gIs��zO����KH�9�SYv�]
K�*�%������Q�����.�9	N͓F�O�2���Y�/DA���xA��?�W�h�z�vC.~��î|){�����=@s/Ic�_a�k�#'̐U����y7�	�qG��u�g%]Js�o�u]M�KWã�O��H�F9��>Z�S�3��[���ӻ����Џ��߂m��g+7;/�t]у�&�|g��%}
&����p.����%"M<��/�\aÍ�Y��w-�E(�-d�y1�?��Df��T�ݖð��r��zo(p|lL z� ɘ�p�H��q�{
�]KDG�[3���:	i�������y�3��4�`�Es����l}E�+,�E	;�t�UXs3Չi��6� t9�����}JV(�70J��H�%��cп�5�������,K��R9>��5إ�Zw;�������Gcʊh��Q��aK,�����}��!b��y��[��t
K�S�Ϭ]��fv��"?��y/�4 �'���)ԚU]PL���GY}��'�1G�6��4���]���a���nqfE��ҁ�N��Ж���Pc�u�kV�<�o�ތ٦ȶfKX�=�� ;|~5Y�����Z�f((����)U�Kv,Jy���
[&�HH.(��f�����sQ���+����Ӡ���:>����~ʱ�p��w�Z�ZCL0TP3Ǐ��aIv��.O�k��/K�L2�pJy�h� ��{�xfZ�0�~���Ҩ;�ulQB� 83���C(j1h����������ŀXi��
XN�:\0����#5�YKJ��	�/gT�ei��kܵ'!K8�u�W�>5i�*�vF�Sk��]��E�Yin���#Êc��]1� l�UB=��f;�pj�3��Z3��2��s{^��f��)��[�u�R�������Ҿ���o�˰q��bi���.ᩫ ]`�hwG^9�
h���l�k�՞	1aߟ#Z�����ƈ��Q�"r60Dj�h��������ƫ��g�_�
��伷��)�+�"{��ʲ��Xz�H�:���K��%gp�̴8	�1l'9�	+���؇�\�D[}g������qC�B���ʰ��QQ=��g5\�kJ�U$�l��Y��ɞ>EN�fGN�ɥ��������	��H�:0�q}H���X�#O)8q�p��\D�6-��%�ˑ.d5*ϕg�k��9��^�qZ���l�M��(��|�ޗ̈́�ds^�(�w������I���β��/P��=���(���(�9u�B�����Te�)�b`U�nF,e!��zw�����qm�^�x$�f��0d����%)p�
~[�, �sR'�\-�����喉0j���B�ɡT����;����jH�o�Лah�i�ӘH
��.�®>tֿ����x���J�w]��B�b"p�Śz� S�gAO���E�L�3v�Z8�f�\[صwSW��¯�C��R��?ɒ�e��A�������O�m��V��������}�7�k�4�}�) �G�ּ�_��l�`,[7�EQ띎���*��e���A��Z���[���|!=�ͻ U|z�l%cpQ���^\�;�E���Mo�+�Ŭ�-�z-˒So���dܴ��4=��� >�D�y����@sc,�aQM�Z:�?��R�r���S����xud�,�ds!�G�+8��
�
i��9��P��'Gzn�P�u�j6G�AC�2#�?:W|�'��+�����T�m�J:��w�J��U��Ĩ{(C��5�J}�h�x`X:IP���2�%��2T���} `��;8��� +l%���I5(|����2n(�����CE�(��9����J���N$BoU�?96�~�U�4i�l`/*z84S��}�.�m]	�zX��^|ex��^�D07�c��3�II�[I�n�8�O��^�>*�]���#Td���?���XDg��7���4�j�S��1��*g��i �