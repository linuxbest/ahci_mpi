XlxV64EB    fa00    2d400H%�_��P:p���F{�-6va��3f|���s؁v���7.�|CU<�6��XD���Vc�8��(whQ��	Wų���|�l�O�C�z8�J�jLbs�l��bzD2��ؠ�.}�8��W���<�ٛw܅ZS�ȑ�ŪhK��? 7(�7�����u�w��Y&�\�����|�\�YW#����s��xT�k���%G��h;ڝ�}�z�*_�tɺ����1ՠ,�c�,mvq?�+��2��Va}�S�Cd�ZRf��_�A8�\@���rfl��p�;r���+#�gl �\��S��� ��C�6�
�,S!5ٔĈ���-�ә�&��Z��&�T��8�'cJ��k��,y�V�1���� 1���qL������@z�oZ{�"*MY1�J�O��V�x�^�KU,W��?;����e)8l)c;Vb�D/cB����,���k���7�J�=V�#��i�:wD�t�L���R���3�!�K7�z�������Jbʝ���2�)i�˶jW�hNj^b+`�3F�0#��(���7�������X�^0�E~�O�����="��dD|�Z�l����V�<��gZ���抺[�v�Y^�ᱸ�X�;�h�ח;T.�\�����`h X�P��dq/�_�ד\|ˠY�j~z�V]T>�%����c�i�.����b{d�Θ����IQ�+	o�U��&F_S}4�Jjh|Q%܉����*��1�m&�A9�b�B.���py�|��)-���a��������vZ����\���v��u�[�������>2^�7���^rT��WF���\Վ�!U�n�Q�x5m�TXTÅ�Y�-At|tu��Oӧ����B*�WȬ��O�/X�9��zj ��j2fx�
*�OQF?7#�a��N�Sof�׹B���v��gN��6���"�4�LK�>�s����)\;¼&n�X��ǳ�:W�zo
��皤�̤��l�0�"M��ē��Q��(f�����)
�4��t�x�G��=@�����~��+z5��>�&AE)�Js�c���4�4��0?#!�8S�W(ld�2�����O,���x��oOXS��'�JMX��*���D�=#����s��"�AE�?Y}%����~T?�>���)�~cp5��]B�S�%!�?�>eU3��ks/�$�6��c�e�	.qE����9p���鸹��9�RCÚ�g"��YW� �NrQ�Z4����\���C~!Y3|T�����@�x���1��yY�>���}W�����˫7�H��	��k���Kv�]��y�j�i�@Q��aka�4.��<�C���w��PV/�$��MD"�N}S���p����I�������1����@�LA�-Q��_�d���`�R��t}lK�;��*�~8z���M�oRȆi�v����w�*�LD]�u�����ptN�"�0<��U�F��l���Of/����yO�P8��#�5Y)�|U�K�U
�/���I�|w9�y�ޡ~Wh�G�-r��9����Z7m�=ƓR}n{`^I��+^T��f:�	�����T�=�ڵ)ǃB2�����=xj޼��=���U��DJ0{ߎ&D��7��L���͉A۵��`��*5�$�m\NwU^��\��������h�	��~� ,	"?��.*8����z�##�@y���<U%#63��N\��	��w"��?�|h�8+�kB�J"���z<hV+�`ꊬ~
�0D��C�ls�P��s����Y߮9�LG��/��6Wbs�L������\��ͥE �_��0w��K�j�ߚ��|4�(q'^�O
\��Y���;��G���)���� �9�I�4A+a�I���@?e�E����G���6gx���4fbpB�D��)TV�n�8�w����)�s�Ѫ��¼��
0I���S��Ņ�n���L�W�ͳ�y#\� ����DC���r��9b�����@�x�U��'d��9v�����1_�*T�4�P#��A3��w���a�-�J�U���^�K��q��@�C��4HǓp��s�:��/�u������\���CW�,o�0dQ�x/�D�%�5�'V�\���nE(�Nо�a����w|�;H.M��ì+BS�{�ai�ݔ�v�m0b�fY��T����h�ʉ�?�+4�L��Hg�Z�ݹb�6�MH�>�v%��Ӑ�0[�j"B#<���;m��CFQ��4���M3�`I�$#��*[�l�!���QlL|����
��
����M�m��E�<�,5c���CD�Fgl�LњC{�[��EQ��s��LʯMj��U�$^}�S��U�z��.i��2?�8X2{�~����-zcԦ~e�-�t)����/���k�uO�	�2���iL�4�������P�[���	��G���z�d/?�G�C2�g!c�c ��E;�q�����_������]�0k��w;|ez���b�g�Gܒs�ל�r=+y17��#d�Ӄ�����AxI�x@��5Ma�ՉSXyh��z���G���65�\7�-�a��ǤʴUH觡f���+;y_�(�Ў���^P��{�F͈�5`�h/��D�hy6�ϼ?G@gjA��o
~Ů`r1���b�ۊi���Y�L!J=��HE�T��^�C��{����V�ώ��[���nyY��ˠ���&��B���Ȼ3MCv�x\���n��q��	�g	K��Ȼ�JK}%+��X�������_�R�=�=�l6���l��P�?'I���4��FZ��s�f����]��t}4/���+��@l���>�g덯�1̰��7>�ܿ�����^�A+�~0Z�\Y�'����6�y��N�=:�ʽ�@���O]]�����<��T�#aN�0%(�c��|N��δT'2L9����R��Hq�bc�C��1wFF|�|ژj����H�C�͵_��[a���(���)V���/��EA�ȁ��S���^q��Yߓ~ {P~T�2k�������Z4�,���ǃ-p��Zu�6�:SW��2F\Aigw��>V-Q6��Hz{��
���Vʷܷ��<�x��ԛY�â��]i��nFk�
����� �*>+ih�ݼ��ŻBs��2�8�!�������Iq�H_A���p0Diy�I����,�d��Kf���;�`����8!ƴ%{���B@����m}���rO6M�E��O�leůCT��p��}�5��g����Tl=����a�F7d�R,� ��{���*��Ҕ8G;��s��LV�t�jx��!���]�tA2V�x�3%�az�t�$o�A�.����k�N������ߍ���w�Y�UN�9�%�0�@����T��s���%(N�HH	g���� �X�y�:k�^���w@��?����g����nM�n3i	|��g�\S���clp�j˨�K�Xjw͛K��N����J���n�~d_Zzl:��'�1�ղ���@��n���C53�I��z�Eq��՞��X�h6.�����̜;6٣��V��5�� b،��-�j��6�ѹ�`�4b�n�=�!$�~��5Km������L�\��_D���ݠ�Ϝ�sL�*�6C6R�.Ξ1��)�S{p2��%�����h��Sx���@V�`Q%�_�阅�GZ��բ6P�>�N����"�8�GTO�ꆤJ{YCwa���AP5��n��p��O��4A!+�>�3��!4�8�*5؞Z��d:v7�O���)���M�	����a��%[<*I�V'؞Ri������i���ѯ�gr>%}�b��Z������x,Ҡa�r,d�7 �6QV V[J����ek�3؅��v=1����D�xJ&5��
EV�<f<?C�Y�q�,ګ�Q��t��SB�<+h}�>S�#2�^��}~�k�Ϻm!� ,J?�Ö�6Y�(�������W�q��.5} "O��WvF(�e/hI�ǚ(_|����A���o�	Nb
mVS'?��Ń�}�[%�?��3���'��?&/P2,_b��JWl�&*��S8:�7iB�%uo�$ߡ��������3�8��=~?�b+�ќ7c�(���w�m"�����<���)|���e���L�'�IGń3�����0�2�hp���UJlF�ӧ�Z��YU�&
�΀e���H�<E7�Y�|�v�D���B�ZXW�f-��SnU\<���8��a:�����9+��z5�W
��i��tU�C��w����!���c�i�ٔ��.��>oH��~�iJ���"[�J���ދ4�bY>*2�1U"-o�-\��R�� $A�ܱed��dP�c|_�tȧ�//)2��j4'l%<Qu��=ʿ4 O�^�]��)���rb�)�
��tG������@�r3OA-C�]���k�����>
f��},V�"�R�y�M��k��N���/����P���N�e
L�Aԧ��>������\� �R�m�SE�H0��2��m��G˪~�a=�Z�[�I�|w'AOM,ĚH��ĩ��Ck�F�XF�C���B/ź`	*�`W.�"AZ�K��ϐ7���5j�ь
VQ9�	%�7���U���+�-��A8&˞硧Ȟ�����	�*��H�Ss����!,�/i�$����s��t�((Z�}Y�X�\M̦�bz������d�l���X�q��	�X����tE�k>I��������V�,^�O�t<?�Ν��F�	�&�VoQ3{,JUԠk�{f���r-N��҈0f�}'�km7#l��ܬO"�?�lͅ�T��ԥc �w�@��f��Z���Qw��+� ����Q�V��������|*ɬ�V�6�^�P��i�Z��������&��)l��
:Dr�8:S�Jx�p����ʬ�1�w�X8����%"�rX�N��ږ���z��]NX�S����በ�$W!kE�L���_���K��ٓw_��	�8�%�	1��@;�n��.���蠶��e�|i��0� �)ERW��\y8��@s� ,��� �I���3�N
���{O�l!������Q�D�(��5{��6Q����}B������x�������r�X�h��mT�~�R�a!IJ�#��_i�g��BɹY����Z=]K2X��w�����e�%J1*T�>*�����B�?�����;Ėѕ��e�ɶ��/�٢�nW�)`:D�$H�����I*�(�n��h�������c���H�Z�6�;
�P��I���Ϙw���<U31�b1|�氈$?M �@�1�/����<}���1-;�\%sN�T;�����Dέ�~4d��@�@�޿�1��V�:�˒�����h��/-L's[���b`[|���,�#5�%o;��7�l��[me/s�����4�"O%�2�$_ʃ�Wgb��o��8}0n?�y��[�n � �D���y�DH|���`үe��^5�r�l$+M\hgE�td.�o���y�	�rb2\6C�C�e�����cu1�T�(C@!�D4�ǌ�bl�����Y����������8����J>���n�# ��u6gX�jäG�^��.�Ĥ�!�7p�(f�#�|j���ܳqh��"}�g�X��t�6T��n!�	����V/��vOP��\#_���'�5��8��l��͙�νz�`��54�^z�{�A�1�6��;��hG�f�^�aF+k��	<t��_ƃ�I�T�7�'���ʽ�2���~�+���i�!d֊�/++��;�Yg͟�����VsY�j�y�$!�%��{��cN8'AXUըjo���O�S���i_L�9�	�s^��D*�� �d"ŷ�G�'��[�,`���e���NA��!5�Wvģ%��UV�ԯ���4���ȩ�s_� ���[��)Q����W��)pxB�N@�J��eT�7�ꦕd=�0�Ɓ�4�m���C���1�ԛ��p��i�x�<�GD�q�$�	�����o��{�T�.� �8�����:G1،|r�x=�5��؉��N]k���M�oԍ;/�ƍ� tZ��y����})�*i����qX���N�ZŨ�4���F-��ɷ(�Q@ͣ�&�`�w����Z�s�@�k���v����s^�Lد F�.��ߌr�̪��s7Y�D\�b1��g�*�Y|X(�E[�]9�LgC7�3����}+�z��5�/������|'l��L�8i_)Q�I�t�����������D��{�9�E�tߖǤC|�ERu���:r_��W�X�x�r,�nT쌋IW��-NI���{~�o�~O�j��a>���ˠ�kA'ꗯ.��U�HNg�K����"��Z��
�{��3W��Gy�Eps�-H���¨�s���=j����8�U�]�:�/_GV��ڋ����Z(�?��=�Q�~�f��(�uJ�{C��S/���ݥ�lf� ���8�Jf�7��y�y�*;Đ8�*��~��rcs��`�>3�U��7}���6�I�F��:)�i�u���"�Q.�~�4q�Hʖg��Jۜ2��	N�7�E�Q��8������zjI#�74� c�X"J�@Q���`�}NZ��3k�����l�ڔQ�����^)�r��Tj$��.~'����;�;P��y�Q���,%[��m��þ� ���ϒF���Ǳn���+�r�HT�f*�ãd.���l^[i;UF�ޏ�yf RG����uOj���>2d�hɜ��K5Na����w"y�<W��N3��1\��v��t=�ŀd��7�5 x��Z6U�b*�\�t���,��z�x[��A/�\��r*��]��KH�o>�0zY�W�8*�O��f;�/�x��  ޷]h�SC$
���p�(�	J�W}Ml�1<a��<��U_�8�=#�[
�M-�z��{�(l_C��jS)#ܪ�`���g5$�%��-�H���
*kFj��1��W���p�8�o����I�o�;�(�%{)�+���%/1�o�?�1]��+����3'G���n'��˻IzlK�1D#r����d��$O�-K�P}�ځ�
ј%W���P���f/��;!X6Rƙz���@��R�j!��7_�����]i�QQ�!���3;Ȝ�A���]BfWB#�ޗ�Eb�����)~Ҵ�#���<���+P��:�pf��X�w��b��
�d3n�#o<��|�9�~�ҭ�52��PI*��/��T��n���O!�8�M�Q��1��L�y_�Y���?yZ�h����X��� ��6��]� v5:~�X�p��F���}O�Ϣ0J����g~��2�Ҷz�o��R��K�	W�&g��W1.`�>`_6��ÆB>�Py�ߍ�y���4[�l��OӘDI��Yp5�'?`|��t�wD��z�����R�º�WpU4�U�?��R�:�F�l�̎�_��b���7
/l�P��v�!��ǥ����!�a�l~Q|�$��(��3�O����o�-�ڢ�=�I>��]/r|V�0��OU��Q�
�)b�#Ǚ^�-�yEǪ^��WBT��ˋ�3A��������N-H�%���c�f����,�
ў��ߟ�����)ʥ 7���ߍ�G~����:�a�"pM2����\#L�ϟf`�h|���1�kn��9vO�Wϲ��C=�
�<��q���[�rG^��� m����Pe�� ��HS>'P�y����z���xrz1�5 Gz�?��ì���O�O���mf�� k�(��2O�3~X
��1�R%��VP��TC�����k@����\�#�� �RH�6CN�0*���MF}���V�/��=�gHؠ`j+�����"N�[�9	�΅�� ���+���s��˿_�~J�BWφ=��tW� ����C+�J�P���K"����p���3��6%+�->��C�
y+�ȴd9��[ʜCP���)''�����B����&�ý|z�:��a�g����EM����t�=C�TEb#��Mu檝a�H3U�B
�W�����!y��x^���
��D6�Ԉ��+��Fiձ=�:K̘��$u����!`y��n��B���A�!H������𵔎}B�楧����D�+��kR�Y��F'����Bf6���MH��/a�$ndw V�Z j�+��O8Z�6�0���rWŔ�	���(E�Ď�63(�@��,��XB�ؚ����$��/oCр�jq����b�n9���w��*�r�Q�c�~��~\ov����ۧ�G�^�KpHDf/��hz�w���0J*���;�W^��2�eCE-�٩�нm	�w�{�l�x�;z��O�x�Δ�<s�����p�z���8����X .T�dmAi��F[�\����}B����\<�4�����sG�_ ��[���8����ÊP�7vQ}am7'�a�Es���9cT�\j�u�^����4�������d-��ؾW7��ⱃ����m������Qp/��@�^5�>Ė�f�H�f~U6~-a8SF��X�+�O�R:�%�m������e���b��"�7h^�%���/�>���Ι޿a�O�c�Ӧ�u��#��/�ؘ��e�i�!赞5?s�l�U�I7�
�~>!H�ᤥU��C��Ȭ�b�w�S�p�9�lLB닔Z��WT3�HU�3"�eT��\�c>�%�C12�&�Z]͗I��K)2"Lh��gf>f����HIL����>�
0���H���Y���ౝ1���yjmk]�,[�q����D��� Ts��!gt�����1��B�}�.yO�`[M;=>�q+�,�{|�;��]����f0�'�Qîc�q����1_+8Z��e�rPؠ�C���h���O=2A����eE�j�B��J�Lp��B'	$^v��=�'Z*C�E�<��k쮅rwKin�j	��죡�JU�w*Ȓ����Ho=_7��3�	�Σ�!<8���%�4Վ��M-��cnuU[��!*�`��*J��<�GF:d�R�na��$�����Z3@*m�H�����@:���2�w�Յ�������%: ���
/sL;���c<���K������ߕ]���ȧA�H���ku��0[��3RϏ5
 jV����e{^Ԃ�V��sa�������|�{��ܻ�OrV�fcx��#q���,a<N��%iˇ���$�Eg���
�v�>��	r��I\w���t��hv#������� ˖,=�[��6Z�S���ʙz�^IB�@І�`j9}��p�7b���|d�&	o��[��	r\M���h"�.���i�;AH=/��-� A�߯��1���c*�dڿ���c��N���̰1,b��t����6�׉[��Lt�ے����x.�B3��61��<e������Mw�X :ļr�$8	D,Hp _U;�+so��<ЮC1W��T3g1�-�����#� ��}��+�e�|%��Zp�w��#�d�˽�Ub�Ac��rϚSW��~ʉ$���e�z?��Q�U�ƥ�k?�ռO������f��|�z��6<��}�ݞ亮�e�=�y��!��&��TZ�57�������r�Aޝ��)~3��োv[��~�
0��q�/`�w[�͢��Σh�<���6�r�+1�2���V�*����ZN
�l:]��d�6L�	��4�����ΫcM�S�����S��Ă�i|4X�#eǆ|���~�8������[��Y��T�e~P�Y�Ȳ%��2�jH���U�S#��
��.��*�\�Y�jz0.�Ӗ�ˠ0��g�@H�KQ��a�m:�Wx�Gr�����cԘ�Cr�鼪�<��\c�H����G2��b�-3G�\�5Sv0_��-Ec�=qI'�nT_,��̌�w�F<!E�8�����(�A����7:5�K�f�V�
�I�:�d����d �
)n���ޯ�I�E%�8�	\�xn��p��t]���-#�����f6$;4�=9r�y���8���̺[��+i3�9W��H0Y����ѭܱ�#����0�J�BG��E�#�nқ���B�JR%%5CS.�7L�?F(����Z�"�M�x\�m9�O;��	��[n���i�/x�s�Q"kT�~�Og�Tm���8+���l؅9�K��s��^��=�9�g3B��qY����K���"�MfR(�Y|,X��i�3ڈڞ�,�����=u�a9���Ǽzd�"�V�^�}�1ɨ���}��z�ۨbS�c���Ѷ l�-�g�ܗc�;�����38�K�.C��4c���z՝�|�E��� ���`���`LY�~�w��`�P��!�աZ!���r�a����ץJ�]3�t��8�T5~��2e��ʅ�^*���9�V��!��tϵ)$AG�%�_
7�����/�GP�c��H6ђ�?�^�y�h�	��{�Z�&3�����,N0�ͧ|Q�LcU�a�ң.rv
��}=Sa+�!�sL
Ucr�R{���m����pۣ ޯF]|�f��ΐ8DJ��P(�����FG
�I?һ;N�)[1�չ����{�G7�	+:	�I$0մ=��(�\3��
f/���O�^���Q	g�\XͩS�j	Yc��U���io�n9��^�i�]4���sZ�/��Wt��K���ⶉ֊����v�*��s�d:PW�$�z�4g�ޙW#�������6�� Vn}+R�L��׼��8�:��������@ϳ�~�z�E���sث��h���Mc��=���E5ܴ���� ����b�.�R��������&�ؑћYw��7��A���rG��*2��u�m^(��m��Db�x`�Ŵ*���a׷�9�Q��/^5��ަ��*���"ϑ������pc�)[��`�����9�w�w���Ŀ����k���㶙� �R�)�BV�����zc�Fٔa��ۯ��m�o��S�HK��bpmU���#	2a�eN�o����E�v�oY��H�v���D��N<�0�Vx�C�p��`���MVI+B��=���a��8##B�:��}yk�"(r��T�nz
���qs[9��8���a���U�b���%zžę�jY)I@��Yӥ�?�h�:�o��?��0�h�'�^��Jl�ˡ������[i�x��y�]�s���,���Sԣ_ם�p6��\�����Jдn����Ou�������/x�K�G���:1Fr���،DXg���Qv�+t]�O7��է)���1w6�r��HP�9v��
��|t�&]�1�.N]��C?�iV~K�}ˡ��a�kS�A�XlxV64EB    fa00    2a30�Q*a���K7��GG��\{��+J҄l�Q��4�)/��wb؞��|���w�a�����bO\{N��u��xP
��n���Y-�<�w���ЧEF�����Ȫa$�c���}�Ț���_�02�G�����N��iW4B̤��O�ǧl����m������ibվ`Ê�����s�,*#�%� ��Yu �؊�c(��􋿉Jnh�;2t�4�M����w��Ŀ��T������RTu�
��	y�����oر�"�70o�$,:��J�,C�h��T�����A>vMN���$ZQ�oP�0\�`�K��>uNxEb[G(��X�sq���Lq4�A�*��;̚�����ruO�l +�6)n���2Q��2e�٘��T<s� #�M�+���G^ۆC#i�?��BY9-m�L���peI?��Y�_3XTP��7|�b�q-����za�թ������w�M�Y	��r]�amG z&���F,�Vi2���֫�����
(����N�x�C]芡�!7���}�c����]"�6�I��o�, 7��`M����UQ�o-}9+�{4v����ִ��P�߶�#9�Vт62Wtx��h�1�#�Ni�秽cC��##C?Մ��f�ݞg�.(a�K�!J��THA���"˞}�أ�&�N��A��֗�(!�E�u�'5����߆�)%U�2	�A�w��n�g�Z��\G� Ԅ�h5o�9�&	#�v��N��L���� nT��;�EIH�-tI�;��qml�k|��HjU�ӓ��dڄ΅[�����(n�1�O?�z"�~��LdZˆ�գcl��6��m�^?�����Q�-w3	�q�z-�Fid��]JWe[R�S�3:%h[߭�u�ܣ�s41��`��xs#��me�:�}�O�S�u�_�[�tۙ</���8� %��	z�v�qq� B���L�R�E�Y��>L��t��F��W�e��p/�K���9.�߮O~�|�Ncgm.�d�f��>}ɰZ�+3)[7 �^�Q����Rc'&ua�x�#$ƺ�t�qX )!w�LC%E1/[h�6vD�_�mn$��QW1O8Sδ�Y=���*����i��C9;�M:�Yv�Gw3�5�!�HsHf�[6۴��T��>��ؽ`Y4�>�ȝ�V^Jf��A�鯹2��F3TJq)Aio*���̙Y�x� �ki��~�E�:܉��NP�b�N��S
�
�V�(�F��������y��+1t�1I��.hBQ��W�akm�?u���2���z�*�����+����Wı�3�`�����z���"=�LtN���[���đ"R�{���02x�>��fMS2z�����#RZ�̲��\Pn��J��W���S�mB~^����7qRX��-���Kaݎ� =1��r�ߑ,0kM90��5����֍)���<����!�W5�d$ƻ���rS@��}�j�;ռ�Ls�9U�1Eճ� . AuH.d���5.����W�H�:��?OxäB��	��6h��<z�q�	���⭃�	A�{eS
�-�j�8 �ƍ���ys #���Pށ�����d5Jf����DxI�Z�oG�|q��F]:d��qxT�o/���@]�9�/���h8�<f�Z�zjk����}0Wq��܈�>�7���<+CQ���f���c��� ��B��a:4���M�+[��9� �	N��=�햩isK0+�f��Ӣ��` ��)�j}�U��*�"Ղ#Z��i6�����n�T�LX6�x6�C-�F�)�%Le޻��q��z�)�(w
�(~r~[�8�|"e�X�Ǉ��]cN���X���ŝ��[H�L�Vn	/3�~)e�i^Ǔ㹦J�ZM{�ǵ�O�>���׾|�x�y�=�P-�Ӡ����d�3�~�'�mH �yve^L���Ef"C'�'�aL1_3��H����oL�4�l]�G�9V�j��췟�*$O"�:��ķ��iwrǯ�e$�y�N�v!{=���N'���A�0E_���%{��ޠz��Ngt��K��u��nl9�ׄhq����ଧ�ǉl޽2��V�`\n����޷V��ٶ�e�t�䩹�=�d��w��r"h8Bh��c�����U�a�L탽Vz]U�A�^��e'�r��0�/����+5qf�����a�T�R� 9�01����Ug���>�A��aQ[��^!:��lR�y�`!�}��s��}��͘ߊZ!piP S�D4��}F���*����HY�_HLWYk�t2��ʼ�Y\���ĺ���q1��g>^���]顢`kV�����,,���Q�:���h|�iw��R�3�J���`5&FY2x��6'�&/, �y�jpx��]��c�%o5P���0&����V����UrI�C����7���RV�
z�*7�vS]�r�),TM�H�	N�2��Ï,=��"����������ǖ�f[�7�wx��kDN�HZ[���]�(��`P�=|X��2^��\��Y�/��y	[���8�l"�S�n�������q��Z+=ч�����D���X����[5�KA� _W̉3����
��E��+�lW��H���+=�ݵa:�ǘ'
���p���$��&ý�Vd�/2-ʮa�23%��l{5�f|0��ԝ�Ӝ���}7�����h���%�b]h�c�U�Fn�ژ�Z��2��Qr�0�����XX����΄��9{M�Ahu~�H&P#�4�N���S�*��YLim����X�&�V&/�p���L���muM9�ٳ���~ų4����OZ��b����t�K�����ל�mR:K�N_�F�O��˖��>���%���$k31�S	��r�d��4���u�g кYm����5;���'��]�K7�|*Olk��KM����?���d2��N��M^�@nn�v7��dS���-ٕ߈S���S��Th��q��� 2����<��j�h��3��䐺����Sb���}�rWk죶��b���V�e�Gȩ�r��©^�D�+k`?���	SqȚO��3���F��F�a�c��يu��Q���J�7����o#g�S�k��PR8Z�ǭ�D��0!V����I���,S�hWvzV�r�s�
1�l窱I��:M@Ny��ykG.;�i{}���x&,6q�mBjVV1B9�r��7�+�A,��N���������k?e0�t4�*'� ��VˋC���Ț���b�`S��(|�N/���D��׊�H�5�������%�DLA҈THt"�������6���ݝ��QKr��>���!������C���aF})�!r+����4��
�Z��p�1�+u�
��K)T~3`c�z�
�k�˚��t>�����`:U�(�u�]:�O�;G��#,�B ��]I��gߋ����@zA�+�f�-L���L�t�o�t��f+u���'��誯Aa�>��u2��K�~{�#�]NS�;{�oiˊÉڴg;��Rsa�J�MFmMu��h�Ɓ��Z�������'naͦ2yΎ<I��%��zcegJ�>��]`O��xb>�8�z_>v�
~�bQ��3��a��/�bI����Nq�Lz�E.0?��ᲩcV��n�
K��ߛ�ζZ	3�؛�	\��0�3��?�﵍	̮���˚ �#��$� ���<��}1ڥ��@�8��9�v�k��`��=�q�ݮ|�9�\3��[S�*0��b�լ B���Z�9O���L,��Sܲ��x�.8�ܧ n�����!3y0̭pa�U��L-�yƉ�a�$a�C�f)�U�o&v�"9��o�<��*D�o�y��^�R�>�4������ا���\ʅj���? �ə�cZ�yy+�!Z.0���*i|�x%=��dm�%7@��+��_U��4y��y����,~4(K�+����1m_����bH�$QV�
�,����k��t�����-���kB�԰�����e�����	SJ$#�0�1��n����7�@`N�<�
?�O�� Kkb�?ќ?O�_^U<)Cc�=*Ѕkn���(y������T�hQ���#p�b�W���Z������j.9)I׬�̢���dW(�?4�j�nIB�?�mK���㭋Y�
ɟ�S��BX����+���.Zغ����I���]�Z{���C��w�,��֧��D�V�qxP�V���F����_��lC���{O�;i�ʞ��{��˃��ħ�Q�q�W2{ͧ D��j}�W�kي4!�6KF���M�du�
��D���+�1��<1������R�G�5�.�7�7�����wd�#8#b�1�sd����ڎ���Y��>�� '��r!R�晕��ǫ�>���ף%bm$�tq� 쌣A��ᙏ�x؍}��߁jt7"�2$����}��"�$�Z_0:Σ#���tPU���01�]�Z+��V\�f^
�B�x�4b����`y/���y��c;#n��y œ+ZE'b��F�I\<��u�����4��6*�?��c'�'\��S5P�w�	�]�[o�*]�^+F2���A\�N�f�Ȣ#�K���O'�u����~�k�M���P3���crl�L�z�J����x�Q�z���t��?mD,�')vk ��V#H����v�vP�z�X��Iw�x�-ѻ�ƈy*8��m�9E��g�BbV��T{�ᰄTZYY�y�W5�nO��
��V|����f ���d�K	�o�K��Q������+-��<t(!�Bz	�Ff��a}��)��R�'�<h� G�����I1�Ҍg+�sz^��h���D�f�.�TD��:
��3�N[n�f.�ڻ3��'j��f���q-ه�4�[�(�ʠ&?A:yH��>�٣��	(4��Ƒ����� n��d��;���F��4�Շz�ˉ>�i�FU��:Ъv�������z�F��d��f\�q*�#�Ax*�[�Z١�_�q�3�-�cSu�ϐ��Q�F����&R\)bp@�S�~�桱?c���9I�[��*����<�2:�|w���
Rm��8*�]l�������q������Ky��gE<�gX��8@?�D��٭ԼL��������e�������	��)�><С���� fe����[���2�2�$���/#ۡP�S顳P�s���=x�U?d�m���3Q�|����aXYB�e�̉�f[
 FRi�>b"ZbR�����鎚҅f���ie�{r��gh3��Z[ߧ'��N��.��B$��?}��}-�	��M�O�c+�s=ҍzm�v�NV������S=�Bz�"�	�j�S?�����XǌqQ�%0e�y��`���������쯯ۭ��!gc��'�����e�J-�`;j>w��W�r������R�_Lۃ��R�2/�B��zA:�զ�l�z�r��� G`)�;�MJ��0��P�Sځ��|��e���lN)ƹ��G���ٛ`E+�%U�#@_
���h���x"�r�����cX��F�����9�Ƹ�k%�Q�;g�¥X���'q���q*�w��1l�|���u4����G���)�����`Nz�
_`�&�^-96��������U#���O���Ʈ��>`���/��r��ZiD�aɐ75̏-i��&%T~����O��L=�<���TW����9N�E��Cޱ�P��_t�f�U�p-��	��>��Ǉds�qu������[�>�A�M�Afޔ���T���h�R��ϗ/�pw�[��f7�	�i"�cS��m�^DRN��2Ì�R#����S_��ر�N�"R��L�
Gd���jEo�lro o���<m�eG�3	����%exo
ђ���#{b���3���_(��=�]o��)o�����9�� (Ʋc����Εs�ǰ��I�}��@���f�EZt.�\�L�Y8��Ν���9���u��)b��`F��37���5O���qK��e�)�����o�(�p��\�Ak�8�t|J��G�zh�t�^�'��F�Qb�lA:����W��#�_3Ai�����!Hw��G�).��\�ϙ�C���c�,Ҷ�^&�j+��sǻw�{|џ���+�[Pp8S���ɌaY=L|6�u����8���0������ɧv���uKW����O�p<����1�� �|X���R,1nj��Ű�n���Znoa�d7�l�\Ő���HzM#�s��Ӏ���Cn.i�p��j"�I^<���)���,6U�y���z��B@�n`Տ������\"<���3�1%�R��Mw7Y}���$�sI���|2�C��2�;����*(v�e�l�Ch>C޷�W�T��~c^��1��iq�!m�x� ����.A�k��Ի�xp�����K&�=�I���A��$�Fm���ݖd�M��ç��z��V�U1�Wb���i�/�� �H
�9�uuۋ8?5i;o�	љwK����5n(ʒߦ��9q�@WB���e�$���h���ޱz��x:�׷5nl,��%�"�����F����fq�u3čҩ�p}*�IX����0�0,���gm�p�Gb�dF��'|*�-�F=�34�xzv�m�*�0ŶX���x�_��/��Gu�i�I�{;v�Ã߮��.n73��F���ɋ�m]�Ӡ-�Bى�G���nC$��Q�2�>v]���ݡ3[�uR˸�`���Q�JQԎ�T�y�F*>]�����ʺ��_�<�����'I�-�@�F�@�!�N��.A��"5�Q�����a٨	@�Ml��/�?h��Wa�����n�����3�r��jOg��z�Nޭ��D�c��Vz˄�x��|Al�9yx7�[���ZҪ�I!��ݙ�������E��+����^�����ƒ42>��='7�j�%�R��\g���r����S���F]e�~GG�rBy��:9�Լ�������8���!���,�C8���*�4z7fA��c&��(�	�'�#���v�o<�������Bّn�A
�$��K;���鰦�
)*?�x�\/8�9�θzN�u��`zs4��0U�)���q(��ςW꿩���TGS�����֨�ς�3dyFg�����7F��0 ��f8�AW��0&P`G2����y���RFt�'Ԛky8�]�W'�hDRu6�>>���)�����.�H�*���~b���!���� ���p(�֜�?�X�����%�]K�-Ù)HX��LA��/u<�(s��Fq�ʅe��-AY"��-q�j|����D���t䥠��ά8 %�U/K�Y�?(�t��r����2XSd���!N3y@��>بe	a �!,��Z	�t�����>F "��Y.�Uu�Q3_�#t9�{v ���l!E�[Qַ@�K1�~I��%D҈i0�v�I�ab4�i�~:X��X��FB��jѦ!���[�d)\x2��S�q�wQ�7�#Q�آC,T�^�2�~r�ěD��p�1�U�M�`��j%�Jv�'��(�$}�3q�<u�!�΂����,b}&��[�&d�tN|=�	*1]�B����1�z�f�.�R�q$�vVwܬ{X���ّV��!�I]VA�R�"�[񘓂f��3[!]�_D�jVHx��˔̗a_6 W��2z@�����82ϝ��}��j�;p����"�'���$����RdЯ�Q�3��q3.�o��/�PWԪ:�"u�/��|�Ec��?� ׮8ʳSs�f	���,�A��ԩ��]�`�׮A7��L�;��U�ʺ��3M���PF.h<��P#O��G0��^�p��'f�[�f#/��(Yφ�]�~bl�ۣi��A0#i"�7j'�@dޓ������V��6��r�d���n �tI��Ӓ��45=E�#KMД=4��m�~�g��)̗h��'JH�m�R� =Z�ηA�KN��G�y~_>~�MQ��|b�����@<���k}U����!n�9OYGP�.m��+���o"��N�M�E�o@�	C�j�mly+V��00��6&�F�f"x��Z��T�i>S�j��2�lew�7?qw>+j;[K� ���+��׳}�j�0����oz����?X\$D��;�0�)��Y��4�?{1�6:Q�ahF>�[t���,7�`������u1C��΃��țCߋ�@Β��a<�Cak��4�C�'�������>���6�4���u��3L�@!2sp��5�;��j�����.���4y� /\��*��[�#�����h.`�Ę�Ӏ��f�f�ԧ�iKD��- �,��o��N>��Q@�Ok���qˣf)�4^�?�.�ǖy/�3��x5��@����i�X�f<�`xa�����QY�y���.k�̎W��X�-��״PZ�+��f��YƜ���b쾜jB�_��������C��C�ǃe��_��Rl���4q�	7ĸ�X|��;�O�x��S�@��al�aDl ��s���Z ũFT��9��z��#�c�_U���_wܒ�x�U��.�:7y������,Ud��d�v-D�~!�B�{9�0vyd�<pNG�xibX<�ъ7r%���1;�9jª�쓜�q{ڳAg�m)\n���Fgf��I�Z����m�$L�\t2q�q���R��q���8JS~o�1���MI������l)SE ��q�6��l�f;o�i O'��6Y�9@��3��,^�Ɓu���ֳ%��h,3Њ�B�x	(���a�:VJ�'�b����v�N�	±~le�o��wP��y�irB���d�d�ȑ3Z�+0��BA(6=�.�A�8|���X��E�w�
�x1v�i�a��2Kmt�̃���؅����.�!��	���%ŗ���=Ի�2g#�\�0�5D^�b}gj���M�rO���(l5O�䋄��ÏW��m.z
��\I_�ة.y�%K(h˽!��jDc��<�Do" ���C�G�2%I|�:��0P��ΚP��3�����*#�C�a�o��������K*�|�&� �$ɤH��)?�u���|
��猈3v����
�i.;�Oo[n��ω��ae1*�m��d��K��`�Li�I;e�p�%�0��)[H_f�����&P7u����f�Z�1�Խd}	�-�kV�=ʝ}rW&e"z\��)c2�v>34�%fJ�EP��0�x���Z��S�zib�ɞ�4�*l���Q�V9{�=�A�D��G��R�d��"<[��n�T�ImݍE"p�&�2W<=T���Ğ0���^�]ys��h�lx�$���N�Pn��#���!�[����g�}�zs�����V��]��'�R[��M��(�����F�4!�6S�*�S�2㽯����pZ5�nl�KixF�'HP�S�\}34�c��8�+�ֻra�	 1���DA�*���fZ��X<A�a�_t�R��]�ZZV���/L�3�{OU)ص�4�m�V�LZΆK�{�A2 �L�ϟ���2�5�Q��(3��|���%I�oZ�fْ�"���m�JH��c���_�Č���ݟIGII������
c�r�6q
�8����V�aFL�19ҳ�2,�v��΀ڃ�cL�T!7���ch��s���i^�M�UBd:��91�D�ya��?\�D�~��]״u��&�,!ΩY��:$�N�������)E��FJ��O�"��m��g�o��jB��V+#�6�yۢ��#�?�u�SP�E�[4Q3o�z"\����uy�3U����˴��n�[2�X�-`���ҫ	�oE��T@9��o�}�䔓�'w�,�����ͭ*I�F�m�s�8\��I�o5���eK.�)>i/��o	��<�����
�U���؛+{��4߽�ˋ<.�LPX'6!R{�$^K���sA�:���GRY�sS|tGV6���S��Ԕ�J<5��WS��s�#۴�X����L�5�hv�aiC�z	d\l��'�7���us���"���:�k�x��Y\6p������C�gD/�Q=�~\���-��P�1]�ٜ�pChT�6L��¦�r��z�H����G���|>ТƼDS�{�'��!�k#�ׇ�I�_p���Re+����K�(�s��7q�h}���r���tRz[h�^���VwM��!��ɉ����CR��}�mbflg�c����A� ��]�W���3���P+N&���>3K��σS�ݧ���dh��tt�@_W6m���#���������R�}��v	���V����r4�l�Z�Wy�t`^g��?O�ʜ	,.��R�z@��"���p�'\�8j�����ߢ>�OFL �JNG�x�!�������~G$5tWI��0֣�����t���Q����ՠ討���ӕ�B�ĊllB�
4@pMU�tw�+�?z�=���)��EldA�;$Xf�/�ِ}�^�HQ�j�=X�s�u
P�P���UVS�.��@��qМ���\>��읏�	\���� 5���2�����-�=�/ ����\�|����M��2�ms	���~XlxV64EB    6058    1320{��Y=j�1���@�g��O�ا�		)��nJٲ�$0@1ƾ�NRX7P���o�aC��.���:&�ZI���
�w����s7A�v>z)Q�5HzK̈́eȽR�%�w��9�E��;Z��̓�E9�}���5]��nx�A�؎�&�c���i���"i�H��ߘ�yʎ�S��wW�À�o>��V���!�ne�`&<���$Һ�=u<G�c��0oF&F�YT���L��Ғ�As���Ǵa�̋is�Sux}tPⷔ&�l�y�ќ�,v
��G��B���:��eV�"��.���[+���0�Z,���Z|��D�3)sg�@�qG�i��[�S��^�(����2�rK��K	~5n���~��BY�S�s̘T� 2��U��=	n6gy�<�?3zq	:�:�$�&c9���D\ј��b�D�*�Y�T`�����$��I�hS��>B���~���)'p=�c:X�?�Hh����}�'�Ðy���jMh<+�����{74X�MҠiI0�g�<����%�X5Y$�ؕS݌��7�J����j0,�>�Q��۴;G������-��B�ƈi�+��)v�m�2��Q�tov!�\�6U�>+���j_�V�R�/X�L}�ؠRVJ��Hb���W�'�����,P�. ��U��67���aq1��wE���)ET0�{���6ӌ�_=�=y�A�k�Ez�s�V#Ua9xoI�æ�Զc"�im�.�3�&?"�i�����~m������򣠔�C�y�b9j8��BF&������lAZ�G���@����7��ƭjz��-��Ct�Cǈ/ʲ�Ԗ�o3ͼ�M�	m���d��j�`5|T�r�Mʇ�R5���(-��ѡ���Fn38k]�R��	A!S�q�'1r�>j|�^,��U���Wb�k)%K�H~&ҁ�)
�m
�U���������:Q�V?��Z�Y���K��>��pv�LI�(!�b����7���ch�.J���Vri�f����� �B�屽�E��2FRV�Y>>��wp7���X@b�&^En��9-BX�n!�G�X\��׽��w��9G�n{����f�;���s�5�M���{�Y�
��ƒ.ʂA�uD�#R6��D=`aᛈp$�� �G#��-`�f��W"�>��/	����ъ�|hB�N@�k����� ��3�TJ���t�k�ksOx��Fg�0��pO��xY_T�M��ڟ�K�/ٸ �1�M8��ۼ��]�H��u�+V�J��]c�]�}��Yr�����?��t��#�;Q Dl�ГJT�>�-k�p�=�.��6��qN�V�aa���U�s���`H���/ï�sOpV5��f��= ��xM5�+�����f#�T��Q�����[Y�hz/O�%���HIj��q��-_����t֑�0V���^x��b�;��_��	J����P�����LH�gaR�K��V���8�@�5:!G��$:�X�$Kv�ڤT�5��,?_�k�.^�ڈ;�����Z\FN��?����s��XG[�R6��#MP�����
9���|�E�$&�鬠����������0x�O�x(����,�O��%@c��R��&�2�c�����zY8@��R�TgܙbpAn���j@�ӗH�Ѓr�*�e��6�� Wơ�lL���	#Gs(��Io4�/�;-������0z3�b�hm^�־�����r@�=v��9����`z�m�
���K�$	PH� �{����������>H��]�l� ?8߯0�a#��n2e��]��[f-Fթ_��j�Kfl�Gb%��(����	5��j��h��Q^i~�{�T�T{���rE�.�k�f������'}^,[L�i2��� ���JgK(�?�D��-B	�IO�
 q�g��
D�\���w2�� �H�ӆi2ԃ^Kvͳ�#��7L�O�X:��>��תI"+o�
�pF/��+2��H�p��Q����\ݘ��ϫ�xr��k1�{��V��Ůj�^��Gi�JN�c�<��d�����Z��[L(��㡺H��[�o	
md'#S�. s>罱0��e]�^i��2ܮtP���L��Н3@:k���'��^�N@����P鵤�Ѿ�����IKBL�pPx�9ݦ����AR3�`�B��?g��w!zb$7�F{#��!>Fȵ`<�b��3ke�R<�r���T3��S�g�!1�ȹ��q����.��#_gBg������$��u>\�f��]�3u:�?�A���|�gt0��6>t�!�B9l��lUe� �����E�ah�u����l�[���]�����_�q��!�F/�F&��#e�}P�m��2�pM:OTW�kh��Q��A�ۡ��2�6J�o����Cs����㻖ೀ�((�Z�\M�0��yL�g��\�m�ُcǋF���C���zy.b`Fr�$#�
@�HM3I\������g_�[#li�gQ�s-l;^�m�s]��m�\0@]��+(!��j��\2[�;bf��1
�(��-�)�0����c{�=�N2�a���� ��B��l
��CJ�Ly�pԃ�oT1_o���7���yW� �S�!;���L�+:e
�$y��£`���L�C(�6� �SfҀ�_��DJh�\��x��d�B�!6�XѪ�Z��.C��]�J�r�R����':��+��ڊG���D��!ϲ�~��C"�&uvVݺ�(܆
l(����}&�}�f�3#���]� X��G(��1xQy�y}ܠ�3SG��x�!�~	�f�W��_�T,з��ZO�4Ւ�U��������Ej߅S�=�Mz]���oB�������u��"�֢���UXi�m�7P�j�p����VYr�4��.)��^=3�]�ЍC�hv�P蔌����k��3��dQ�/��$�!`�+9�y`���%�s����63m��hTk�RAۧ��*P��N�!$�#\���]G57EɄ^�h�-�*A'Acf��#�X�&�����i��h��P�=�¸8K�pz��� �w*C桶3�"����
�?����b�U3j�cR{�zm��PI�^�����I�+�u�s�h��28��;�"�!@p�I7'#���/�B�@`�{�9����c�T1��t��%��0
�����/�R&!�_�+�*x��wh�.2�qR�N���s�]��H�4�C��@{���
���lQ y��ng�����k�2�Kl��q�c��B���a�Y^�c���T�)�i`L>����JNIY���M��1�����N�S JK
k�sT"?�Ἣ�&�4�v��O�}a�=��O�3�*5�2����Q�ס³|�����5/�D&2�j��2�Aq@�=
�J��1-u�ppԧ[r&��Wy��ǳǰL����t���k�(+g#�kE�����nC�jrk~�6��L�c��R̺��@����c�p�uw�&^����^������'W
>��!Q�Fx�����"<t�C&W��9�D���(�&V�m��`m���r/���R-��\�L��Ȑ� ��Ҁ�+�kʹ�s��ΐ>yi��-1	�"��L0Ł�`m�ki"�����j�	U�`�p�^뵸�Gٸ�����Ԏ��� ;��Rz�7b�����/w�Ύ���˟�7�k@�:�@�'�f��<9V���iF6ٯ��{9!�������Ǩ����qv s�Iۑ��<�w��&�`z�(s�Wn�ȱz.�M0����A�x3��
 Wi��U2R^���ىv�|�"CT�����d�1� �{��'��P4Z��Kľ������cJ��~Q��V~Y
9���#i��z���=춇��%Ĳ���ͅ9xaM�����h���D,\�J�n�P�g����YJz�@&����~�g��C�����a�J������4���
D���?�'KխI1X;�ˎ��JW�>ͩc��4����Z�Q�Ի�1����8�+���Mr%9�#i���^���n���S[^�&��,��Z�c���E�mjX��!�����X�ӛz<-nHp5��_�<a�D�
�S��df��9^7�%`i�= 8��O��\t|�챀���U~2�����Up:xatv�wp�yt]WC&���B([:-JSҁ \��j����{�>+�(l���d��I?��Q`he�?Yz��C~ZfnLT��#���YK�\I7�;��h2������)�N Uy�8�p��dzM��;$��7��{#8�Ԡ��E%��~X�A|վ�l��%~ U�ur�P8'L�@`�3SX���	UL�ջ"�a8,�Z����&ڑ��>��P�`*M<FV�v�8M|:�[��%]��̕lq��Kf�i��a"�sLL�m���n*�jq�C��%�o��A�|e��v���Z�!)�?	v6 ������*H���y������Z��S��7!G������0������0�i����({����1u#�����Ԉ���e5}��mK�g�]�'k(����'�ȇ�%Qle��{�H�C#r��OVl�����Y!�0�-"�W�;���#˚ ���w�'X��<��s�����r����O9)6	��k{�<)'�I(�9[�-�y���.X�xe<�z"�s�\�g��ZD#e�6�ە[��]T�H��exN�dҢ����i�=ZRC�vpp�PA? s��f~�f�d��10mA
3�F������N������x�������:>La0jK�"�S���Y�}�����d�!���ją�		ϱ��9.7��<l��ۡ�F̞Cfks����I�a