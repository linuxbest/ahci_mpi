XlxV64EB    18cc     8f01(q4ɢ�Z$#�=ʡl���GA�-�e6yg"Y��̣�;� ܭ�e��S���2̪�~C�;��?�.@���8G�������s�Ӄ��y�әc�Z����9��îЫ�Ϗۺ�;zdZ&ߋ�����k}m+k��񟆇-T����9�Y/���g'���dp4z�MF�K�M�Vw��+���,+���K�Qz����]
�rPM��N�&�Ю�b�q� ��{�l۞Rڡ�;�M/K�9�%P�R�N2��8
��i��i���	���xo7,)	}(�yp�'
�-�&��_t����R1ؘ�~k���������ȏY�"�+���Juim�s�ɓA�W�zMqE���w�q�U����=�Y����+�R@��!�;U�PZ����1���):��-�+c�l}f;5N�dI�z=��Ȳ�P�E��W�7��]���+e��9���5�Eo��C��!�V�6O�^}
���/��>�(�����=vwM��م��K����yK&��"j��IX:o���1L:��(��M���q��/��1pkY`	��׏�8����n���r��X9�X�����q��޾U�}���}&��WAgPl�/�kZ��v��
&����`�ν�z<2���3-L,�z���"h��(���I[�y�Ӷ��{��0���Kײ���abQ���:֊�N����0��r����\�/��V�(��/cr�s|�A� ���V&�F�吜ŹPb}��Y��+ю@M�5P�e膧XA��0S�~��/`ޑv[)#������k&۩\񑜿���0��y���ӬNns,�I+�%�
N�+��|0��Ȭ$��|����2P�
�Fz�p4ځ�-�G�k�h6	*�q�����R��H��t[.L��� y�"�Eg8xb%�A�/Ɓ
�F�h��`��@��&1_1a<"<��ֈ��d�&ގ}��$Ӻ9`i��직/� �naM�ݣ�^A��7��H{$Gq��dv�S1l��0ʼo�)���f�jtR~9���]%�@�tG�c�_�}b�N��.�k�s���݈�d��G��
K���-�y�����_�Ns��!�Q�9@�����QZ��^Č�� "�c�^J����զ��G�6e
]i�is|QV6j�������]���=p������kY����̓��S�(�D�A�)8��ӳ/�o�eB{<�$�ib�ceF{��?��]� ��\�tD����ǉ*7H�;��_��lg�0��H��JD�B_ c�HBV9wGw��#V�N/yjn����K=�b����$Z���	�<���M�s�7��VV~u��-`����� ĭ�3�����UnI���?B�L�uF�([��&�xC��W�b��K��v���!�;�vjՈP*w������b*�\-F���'3��3�����:�L�'�ݾ�ƿ�I�.�8�3U��߹�/N�7�1������.��/]��J��������1���{cG��R��U~�a�ZF�M�h�7#��a��>�@rO@�`w�Ȕ�����thp_'G��@l�֝r� �_�;�U���EP��d
�N"N��5����}۴�')�nn��v�ߣH�O?DP�_I�ԧ��y�<�csKw2|"طv��w�d妏A��d�
M2�F�
��|�R�ai;^!pw��Ft�|�-�2/��@� ^��:rq��� �|d�X�S�u�p�~i�B�_��a���Nf��;�b��y��{/4.��l�3f�C�L����x�$��Ϧ�,<2Dg��%���le�����2�m:����҅%�x�{r�L� �Kbĵ�����ۘ8a(�r=�*%��DM{
^z�K���^+\�+���(����獊k*Zʏ9�Z�֪�ۨ4n�$:5Y�M�����S���&L1F��@�=Z�Y�nס��p�5�Qk��c�t���-7����[N+O��x����㪻x��@�I�`��U��ż���8�u���Y#-O.��;+�?	��"LZ%\@�]�~o�����$B0�s�D�o�]�7� �v@I��� �z����.�j�'�k1 ᡦ�k��>��b��p�������eapS��koV���N'U�v1���%4��5"w�2R�vO� �ctl.��m M�ɂ�����I�tc?��r���K]x]J6�����˔Hp�d�_2���Fب�@@�	�R��@�j6g�Ĭ϶�V��R�