XlxV64EB    381b     fb0b��	�`\�=?/8���{�b��ܪq�ܪ���a�J�f���vG	�0��־ 3�Y�j:Ԁ��Ѷ�N���,��5�'������˒'�h�N&�bE&��<P��k�����u\}�}��m��<���GW�R��N��g�V#���]��M�7f���m����4g�؞D��}��P����!r���m�ku{�ha��LvS�������Շ��K�'�}M/����aC䭇=��������Qj��Ny\B{��z��ʁ�g���$3g��#C��֩�I���4�e`�����J�$0��q�����C&�Ky�� �mL�z�>L��&P��S����Uf�M�����.�6$D}B�~�t�ht�������q�A(�͢����r`pcr��c�o��DL,�y�%���ħ4�ac�)C,������n#<[�a���|���,���t��o���3|Z�δ���~�^������YD� H��$;{;U�p�1`�?�@�����+W[!��(�E�O	%��T��D��,&��.��jI� B�1?���Ÿ��q!��1��>dD1/�HdxF>����G��s}���}��s ������ξ�/�I
��`���7�3��h��E�.RШ��N�s�4��"�׸t��u,�����jpr/���si���#ҨI=�V��ꉌ�F��$xx`[��óG���K�>��8�pܹgR�,o�����E4��ߕ�4d�G���k����m�� wx糈08əI+��6�ϱ5�~���2����խ�o�w� .99�< �%�)V�\�װi��V��	�L��Լ'}��n5�z��R�n������5u�2U��@�/�`��.���O�&���`fA�\M|��aU'󋦤�X��UV��t��
�F���C�8霿���?�H>�tw�3�Qu^�l?QQǏR���@A�\b[>MPA֨��v�6��G�PVb�{������s�u��k� W�v�^]E������#~O(�
A���z��ťn�^�W�=���ם�NodX��;��]�k~�Wu���2���n'*o�vߨ\36��)�n�� x.�� ��㪙��BX�K�_�6i����GrU�&x$	�zEj���B�b6�h~a�b�mŴ5�Ʃjx���J&����T8�)W�)5�Z_�ƴ�r>\�bX��8���E���,�E����O�&FiO4 �TMa=���K�`<��~�i<0�EQN��	����$����
�d��¶F���V�V`g�����W�.��ʹ[5_zV�� �+���G&�}0%�Ntj�A��洓�29z���a�$��%Z�L�R�^1)��}��{g4=?��O�'�Xb�E�`b�P��~��wՎG����&R�۝�;�d��̬zT�9r/;7���8+���.�MNX:b�QVB,l�{��	���r���W#�5ԟ]��+��Y�ꇑ)���:����=�H�?�iȨU��I��oVr�H������}a��a�v��0�����C�cR���w
N$Y�)=�r�ۆc �'��9 ��!��:z��f1��M'�"v�n.�/T�y����+b��PXD����1mW����;�P1�V�x
�QKD�gfO!��^�Y^'}&4x�����V;�P��Ml]r�,ad��<�`��i��B�������Y�hHu���4C;a6d�99?�G����� [��ih�3q�h
������1���d��`�^�a9�Z
N]6+)�nw󁍞6���>��%V�|�s����r�C]��J�eZvJ�.ʛ��jw3��ϭ��R�6"o�^�/[�N�۫Q!�O���w#��$�-��D7?k�M5t$f�O]�~�V���,^ʗ ��=����6CyҒ��"0e�}�8o�aF�;j��<dkFMRAL��C��%���2Y��� nEM�DP�#[���:����6��
8/	P������z�3�5��$F��?�9�J�6�V>e�䙍�������'�g&?��?��J��Ր|�YЉ	U�1D̠4��4R�c�8�>�[����Ѝ�5*�0ڰ�h����Ēq=���	V�����^�^���;IV6�0o}=ض�r�U�-����ܗ柔�-�0c�:�|�5c��~q�dNR�O��%w�._U�f3ʷ?KgJa~~�$�9��hS�[?��P�R�Drm��z�Z�)�1�s��m7���z ^��K�Rb�z�%�}�����<4�Z�Bl�̖�ޛѭg�t���1]�>G
���&r9d�������H	%8Y�m�W��e+�=���:��j��cdDK���>[�_�"w���Cˑ+9�<p�R�E�nj�L���	.gE��	�`4����7 ��n�A$:�>EUZӊ�/feѩ�{�Oߣ0
I�a���44	ӵ&��#�s��	���D��d��1��E��uo1��\��r�"�q%8��s�}�œ���"�����o�YJ�G3tjf�w�v�p0�~�߽��Ծ��;����+��"<KV}ۇ�(4�(��z����`X��a�
u�F���vԮ-�U
�~o�yW�%V^5 ��R�}*<�*���ES��֢^.��C��Mr�>7�{T���	�c�\��EW
�䲗��Ւu��N&>C=E�(U��*$�u�X�c�(��LW�缫���S,�:�win����ܢ�F�(Z_ޠ_A���p�uX�R�]흧�]�ڥ:���n�@��y��~��Ժ����G�#�2��B��F�3="�N�:��֋��j3G'#	j6��K��w��{'tQ���h�=�"� (0�t���ҊY���8\���Xu/��ר��_i�L�E�\��m������iʪ��2�z�	d��O�� ;�D=����*��M
�˲[/F�Fc~^�Zp��||�H�O��&�ҒKb���DL�*-�E-Rר��,�MUDa���u�̶hA��Sx�) ������O?�3Q��<T��d?��Z�{�N��H�����&��Z�Ą�������mӭ��#5,=�`��6�l�N�o
Q�:f���ת���!6[HO�͆eԧ�TDtE��z������f��:��R�V�:dn�jC�dbj*,��rf�>(eI9m�Szծ�=��l�=^�_������T�Yv�+���%�`ׯ?7��xrT/�+�#�ע�¡4u�4!�'��0{.����]�ʅ"7�?9|��nz<�;���͛�Q�o�������by�V@+l���X{4'�!L�أ�/iW�ɠ�YuŮlA��E�|8v�Ey|�/ӔL���+ p7�֠Q,�Pq�(�c7ОN��f*!����p<���8������b-P�Z���U��M�R@*���|�����k
�Xc��:��͑Z|�,���,�n�\�O ����r��V��o�8�H<@��K�"���n{:�	�*��t���Ձ�%q���Y-�u�Y��3��Y�F-pw�]��C8�K��׃�K��'���lD�u�x8�Ѧ�]Ζ4�-*���	��T��8Ŕ��P���D�����1����<��1��[��1������uw�i��^���o]��ݾr��N�}̄�N��s���������h;�D���*�h8I4�!`0k��p���3AJ�̵ �yu�&	�Ԃ������\-9�7m��A�5t�R�#E6��0U؏6{���㧋�X�e�^���xnY	��A`���䖻a��H^ٿ�&EQ�P�2��\Ǽ�P�Օ�X� 7� ��GDI��O�Tߖ�Z�'v��
�G��Dk���F�us��P�GFm�2��rr0Km:�`NzQ�b����^���]�t���m[$8��Ҕ�����z�3�;�n�!�9 ^8�*?w�KXŲ$Tđ��G+����=������[#�l%/��K��m�vC@��Q�L̰���d�