XlxV64EB    6324    1730�9��͠bP:��l��^�0�`�y\˩G���}�Uz�k�E����j��`�p��x��Ǘ4�l��;>s�/X�ss��'�[���Mwj��ϐ��R!�
��ܕ�G� ;+P��l��EDx��UlE�7�nH��p<a;����H*�CV�ڥZ �E�x.����HetXdկn� Y�j�3�΀4{lay΋I����%�4N��ƹ%R���n�P�+	���;����6��fI�I��k^+��R�"帅^g�x���M�q~$��®Ԕ�hE��m�'O,s'��Og5��X_ZB��#l���+�^��jB�e��y��#��;�<�"�k��N����8-wБ��$�?�Q��fC.a�Qߚ�����3�������9�"�# ��h��Yn5�N����%�
�S�2'�.��Ďf
�\�\tUV�w7e�لN ��#kK��U����z!�`�jSUc��ۻ�� bE�'��gf��E������$��l�3���h�[貿"�E��0���O��E�0���a����0�c�K�mǰ5�#1�Q8�55y"���p�2ߠ���H:P-^X�N��`$�#p�UV(��C��1����~�C��7jBt���(*ޓ�&(�N��J�5x��-���@��dj/��~���`�#z����g~����_1ȷ�&�E	���p)���(�I���c�@4"@�֩�S>�;�o��8���c_;�Tl�#�]�8�d3
 BZz�\�Y��E��T�kW��SD���I�3���{��0R�P���`�}�����=��S�C�hN.�j|�%ޙc�.���N�u����(��G\dY�"� �XT�Ih��� |dN��Ì��5�e�m�M�!�kh�Q^�}r|��Ը��bX.P�U�Է�u��C�}Z'tP ���TJ�	�\
�ģ��LY7�j���G%^�*x}���38��rӽ0�w�hB�;�M�T��\{���Q��eI�����Ր����IMsY�᥀��9lޗ�����,Ը�Xb_S�<�d��W$6�����3e3��z<���8��dv̌J�BH�Mja��A���
z�|�q�'�xԀ�^EXKihg�Rm�+E@���s2��j��,5Q��A�p�뙚e �l�ZWi�3Qx�N��S[o5���3II���#��&Э�s���S��]ig��Ӧ�h��Aԃ��d E��Ov���kIV7�� M��12��͈���>A�r@�Q����{�]�RuPB-~j�/�A�h|Tr�:����Ǿ�D�վ�|3{E�9�s#q���1T}�tĤ����h�JB���~��Z��5׾V�2�hDy�x3��0A̜���y�\o�" _�Ngɒ��>.N��B�U�^�0fޟ	G8ra��|���°�(�ݷ3S�'�ˌa���P�qe)��t��jؙ�5��d=��Y5�:��P�޸8"�:���Z�}ď����m�Jx7�@<[�ә�`� �ɔ{�xL%��B�p� x�1����c���P���9e���Q9C�F&���f��,�0��P�F�y��xC��F:ox�0,n���}u��F��r�2!y�G� V��$!�v�t��0}��:���}��C/�P|�aYQ�
~���G�� "zL9�|8#��K�j��ё�6�W\+^�5{�R���1���!�j� ���ɼ�޾`�`�����=�S9��ș��"�3�������tA�jo�x}��(����z��=��k�O�mV���#��MWsБ�g��;�2����X�35��oػ�˂���K�t��	H��z���������A���mp��x�=�{�_�岩�@�� � ����+�آq�2Ўz���3��Aj����Vqڪr�W�����IZc�s��R�͎�1m 4��!WDP�X�S1>��G�n�ő�CyԔ�P_{P����n�����NA`2�a�i��7ʡyN��/���(��,��9r>��c�늬SuPBJC��JPo]�]�����nIՖ�X)�8�qI#w�O��a!&m�M�9n-
�$Q��I�P� ��ڳp��פ�ئ�� `ԿT���H�~FH�g�
qu����'��f�fp8���G!E���2����\��(
�m�d�7�G+�>i�o;]7��@�n���Q{��D�Q�1!�{=gG�h��O�.@P����v��Z9���.����_�nw�:�ex ͇(�3y8�!�X�r�;�G6��s|���ߚ��O����%g%+�/��|�ưq���׿�}E������"����-�:��L[7�UI����Y���A1�А#�9����"z�~"7���E!��KB�7�[$��,��J������}�=��*Dt�ɒ��L+�ՙwJ�h��i�pd���W�b�pT�X3gJ8���u�jT��^���{�@��_�l,�t�Mm������x��F�F���;^B������^	�	��l�cC�=�"B����/��5���һ���|�Ck�O�i�]���w=�}��Z���x�4S7b`wu��C6��f30��Y���xj���d�Y�*5�1|\<�9�+�>d��_>��r*�W��8�}���M�7�ыq`̦�fȀVD�a�
wg=�eG��Z�GD/�g~@'̘�Z����B���/�E�D�����s�tvo	���a�H���i�4ѐH2��2wU+��uG�P�+f��
�%���s� �z�
��54$�e�P�V���Y��Ը�o)T����G�]m�1��  �L�rTt�:+'�X�p^���^�S?�Fգ��̅�kz�%nf��kۯ����~�0kS��'���b�����9t�QB�ǰ6�ׁ%'��8^�LsO�*佖e�VM�l]�e�r�-^F.>�����c�
j�e7��n'b��՟fb[����E$�&��d\�]؀�.�3�_���ɛ*�de.��+�� �����-�|�����u���,� �k�6���a��8}��?Pz���g!��o���&��cu�]l,0xi3-v
S�J������ҫ!��$D����e0�*C�f=��l@����ψ�4������\g��u�@t�=��-S��9� ��K��*R��/�.01�p߾�5*۵ˡ�
���	Q#�^����f�+�N�����+C��ݿ���11�H�5�q�����	�s�yL���e��	�H^WR�,:c||��R�J��#��~�M"�Fg�Me��"�����>(��l�E4Q��H-'�:3����6���<#o��m��l���E��ut�g�N������ZM|sNq�M3k�I����Q���CNc���5
@�C�،F"�w�RO�@������<�;�G�Sq�6���nR�(U@���o�q���Y����q��؟��%0]R�6��{�-��!��,��=	'���uf�O ����1�C�-���!�	���%��kݹ��9A��P��c2����e?3N3Q�6�â�iO6s��g�����pa�y?Y7��9�3��'�8�.�9'�g�J�a��]*(=	�I	;'�u�ǆ�սQR�(=�HO�k��� �oW��wR@�4��"Y��Z�����j��\�T��16u�I��«����=
�U?qK�stR����Xݐ�^D���$˞���_���ѓ�i	����N���)��Y�܍W�O��;S���=��+3T�J��xNƥ�?�#w��_�g>���=��I��5�*�⵵t��T��-�꒧4#��Vb���G��o*�z�ي��vB}<��+�\eN=fr��-�Wӯ��]�[(�/̿@�q\�<��}Q�,�lK�1|������)GD��%�j�E:c}ƿ�!�$3(�1�@�Q'3��V��;���4�_���^�<|K�"�M'
C���У�6�քITjD��0������0*��s��J����R[sN�l?Y�&�������	r��"E

�X<R\��dV�D�v8���W�)��m<�8�c��R�����Ђ��S�T2ݤIሦ��a
���F|ʍM�;�h2��W��,�Q����"�2s�כ��?l�B̿hP]�&�4}�-gW�+6�̍`��������1�s#sY.P^g:���s���o�M��a$�}�/�:����]��<1�m(s���aPC5+��(6�FJT�S:(��~��O�${^�%kZ�T,����yV��%'�5$�&�8R5�R�=to14f�b7I�	�H��{&ݔ*Ɵ��|��(V*iI�s|Rx}�����������+��N.k5<�/�Z��Hu@��� �$�T�Q��������o�O�8��B-���x�0@��9ʮ.P��}����N-Pr��$S\>�r�s�n�4�P+��W�*��;+.NP��IRd��Q1�#�Ӝ��_�*2<kEhӷ�n�F ��'��9D��~"!-�4(@����ܢ�X2���qP���+n�}��7-9��} ����s$�}�).��k���*��g`c������D\\+�S��qX����O����o���,����8�%����t~2���_��!6�/g~r����]#��βdZ2N)J�G8\:�y�Mn]�\l������D���>�V@%N��<7J"����8��������N�n*x{�H�~HDg����k��\���������ت���L��%_�]�ҋդ+��)�`EO�',����wx�p���%�E	g[�(�9œ���T�kQ�u�u�S��9�B/I�� ���F2��_�����^�Ո�Cok�ʖ�8/:)���G��0�S��D�(����&�U��Y;���\H�c(R(���gTC�����nVGg���CI@�!_���
8piے��l��}O��HA�@���i-m���g���8�Y:�r&Ex�g荠:�D�?:����0��&��L:Ӱć�I�d��� ʐ��ͪ}�� Ԑ�7�g������A�v� �5��̳Z��3B���+��w�q������Y a�j�[���/�u{����+_!����[�-c�*�V�\�t�B���B|D[\!�c�c�H�ُ%�D�5�遆��/^�v���n?{z=�\�cJ����jb�q�~R��M�]n|."Nf�Q	
�4 ��"�48����LN����~h�o�����k�8CM��w�L��_;�"R�J��\�~��)WK��LJ�.֢����D~܎�R�<)qL!#���[�܋�Q21�k�/��r��&��U�4qd��"���/_u]@�u̐=����+Wf~�Ԏ&+Es�NQ�����4�G��4��Q����Ǿ�vl)u4p~t�����UÉ��s��Y�Z7�eGQ���de�Ӎ�l��Fl�3<'�Qjo�X��D���Y�ʤ�F��
���DJ��$FiP�^�_�p�ش���_����v��;�
1��M2����.�C�9Dv]���Y��N�Զ�7�o�M5�L�4%kc�=, ���ub��>KxB	�ü�w��py�a���pV�ED���񥵕��`�.����d�DX2@P��h#���n�<�7OX���� ����C�#�w�c�@�ŴS��������@/ΥΆW��ԁ�U���<�<�͝U�(p�[��+�F<.����ݖsf�~��ߗѹ����0Cz�����\�{��
'�YZ6m6��"���iL����gh9�倴M�uB��`�#�4�2mA��D��v���j������9��v5�P19�0