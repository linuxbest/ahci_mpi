XlxV64EB    fa00    22c0���W�GTU�����'�V��.���GQ�Z��g1K�[��rcf'5{�����\
� ���u�L�(�`�W����L�\�99�-|��*�e�&�>�w��y5�z	�P���k�ku��'OF��Kg�z2%���z!P�٭��WTs4��W#I	�oᬫ��-���g	��I������X=p�WA℈L�13D�)��B���4����62@�Z=�ǩ������m�N�
#"���{ u^~�����Ρ ����=���.��%]�� ڱK���~@�s:k����JJ�-��ۢ�4}L7���`�̛n��)��ѻA��y�)Pb%������KP|��+��nk|��@bu�3��v�Y�r��=,E���B� 5*c�Hā�p��Ϳz����t>I��K'_�v7��q���f.�"z�qn!!��,���� i� �r���;�~i���,�Z�n���d(���cی
�.ӳ0��[Y8���$iJ:T��5�9�FWw�o��h����F��巟D\��.L'Š���t�H{�Q�`��T?�T��믥��T7�rI�M�{z���m�P3C����q)��<��}s����v9��0��u[��`�YP+����9�(�%�
c��mh�*���~RO�L`�u����na�wn}h��K|��d���G;�96��J{�q��_�Ͽ1���p]I��eX��֓�4TC�q��D�k-)�*0�l���K��%Ǉl0��_�SldtHSh����{:��DƫB���	����3��%L0b�`�����穨	�4���1Pxqy�:jȑ'iʑ� ��@��&*l5g����˹"'��B9X���K��Oe�[Bgy�ٌ�`!��U�c^�kHS8=�&������)9+ˬ����K �q�I��fK	<IV��L�ʪ�(-���2��ɥdOԻP'H�IR��
[+�O>�ܲ��տ,~�M�&\��˾�AFY�iY�n7��Hm&R��L��E$��w\��G�>T� �˼�g��P�c��\�^�O������� ī>}��P�k�u�!�v�0{,��o�@9�������.�L�V���O��Y��~՘�8R�-�%@MJ��/�0��<�^ǂ�7k�L0���ͮ~t=�y���~�9sZ���ߧ��'ѽ0��r�W;"M��n���*�S�t/8�n��E8�ƨ-+C+��t}v��:�9ɘ��`ܵb7r?o��'�=�	idT�����.�2T��}W0�k1u�A^��RDU6��7=e�i������!����e�q+K8>9�v8:ΙK�ꬤ��$^�em,~��O� qa~��<�[�����3���Ud�~�c
,�q�1d\� �11"6�o�F}�|�N7�~,؃Ήl���n�S"�â�/T>0!��L^��)�`�|Et�)y�H�#��4�`�@�6��&����<!2��ѫ�Jss[w��s��4�Z[�9�s���$8�t�l��
���B��P������<�
y`�@\.!�2Bһ��P6˦���������N7 3~���pM�=5��;٭&���rȕ�.�.�L�/|p�៣"8�8��B��r�I��MVd�(ֳ���9���ØA�W����$�
��n(�p������X�F�ힽ7�W�_E�:�w�O<�Bd��v�R��%�1rB����bi���P ���5c&�J��"�Vl�1��z5��G�*K�"p{;�Ρ�@���B����T ���æڙ�r�p���Hp;���d�	�j-�.[�^�mȫ��v�� ]�5��H���;aVS��5�x��nr�<O s�ndg�*�+�Ú���:T*n�����a���O#&~�1'����G'�ɑ���u�a�|>�Y��>X�޸�4�d\I���#�ԑ!���.�~+{y��H�A����/�w���%|��W�A�؅խq@�酨������'��]�:�X��7ﹶ߽�P@��>�w2|�'݆ؽ�/@*`Q�9�Y�@ţ�yD�@��?�OdJ,o~�����*�$�qN��Z�Y��nYx�X�C��H}���b6����
�+cԗJ���c�k����󏌡J���Y?9�������.0N$��pVգ�ՍT�p�Ղ��C����S���RB��ea�J�.�H�'�
]vl��j+��WW�i�����T����������iꐆ����߭�F���K{}3�k�e.�#W#�א(�jE?#��>�f���4m��M��1pB�K5m�o�cP.`<<{�!#|ѝ������C��?�������b`�`����l���u��ߥ,����
 &�:�1��V��SK�'����'�%Ԛ?KKC�{�K@�lt>�ϕ�W��r��y���=�VHP�إPň�ފ2�	g{.���U�]R�w�=�9��*�b�	���y�7���µ�Z�nURl��z�B��hEͅ�t�[�#D�ڍ�f���{i/:ߕWIc|���'�w{�"9S��}e�����^O1������R�'����{ʩ��nИ��A���=;ШH:&5 ���u�2���ҝh��ސעe��{�4_&9"E�U�՘]��:w%�	�%l,S��A��%��D�ɴ,8�4OJ���Z3�����/>���x��F2#�ނ1��c��$h��0@)���%40��&�~�U��Q�Ǚ�c���ہSA��[�`��#$ ��α0Z
s���b��L�̟��*1�B�%�Y�	3Q2����Q�ĥ)�kŹ�wW��V��Ի'�z�+
��J�� Z*G8���Ac�FH���8�a�Dz��2�^,y�OY����7yw��NC�@��i�
��ݝ�r����AC�@8Z���f�m�nu�(��Q����p��Oi�V2��{v����8�����E������[ҳm�A����d�j k ����Є���C�%������!�$�"=����� ��⌫��B���9��.Q���f�h'�J�q����E�
gT�n��`�V��4�W<bv3�����]�t��*k>�cWV"��������i��&q)�4D������b��p�lD���zA�?�)�|�V�i`�������)o'�Z�t/��	XKK����G���h��n�-3�ۍ�̙o*�0��i��Gm p&p���0��錴����x����2���j"7{�!��;(�4׺��B��I����/:y�n�G��V��͊���lU虢 -�GCȗG��z��U��G
n���$�2ﶝkn���<�^#Yb�UlQ�<�*��y:�/-��DVzL�P���ꦷ�u�?��i��|�U=(]j�>r4�쫳��� q��Wտ��Vܻ���m4󕒑MY�lU�N���.��M*?
��������`EB�df�G�����,�-H�U�]�紩V�T�0�F����_( �����c���{����(�v�x#��i�"�SV_�o<�􈇔�e�?�>甡�F�3XU`Xн(9X��Юo!7��]�V#���ULh����H���i�����o�$�|�^�����z霖�O4i�#�:�m�8e��J<WR��\wȽnWG�QU�0��\��6��Y�n��3	 ��BDɸ�Z혓��3>��SP��0�#�z�3w�F�,�눸��Χ�.��i2�: ����f\� ?�cU=���dr���CV"��� v��\E�\��vVKjJ��U�]㝸0���|�r��M}Y!Q3��b�����w�+@�{���h���`�r���U0���eݲ ݢ-�:�rk/����B'�?�T��T@4�X�Ē���9��޽c�O�_ބ+����,�`s"BV��Ȧ���`�q��"��Y�˪M�є���'��!��կ���.D]wp�������x+����)�U%�`~7m�YX��N,
��
z��e�Ѥ��5�Jy��;���\32�p�!,Z�ޔ%�o�o��n/ $D�o�0�;@��|͌> :��iu��U�4G�|�IC����G[=�δ�T��U_@��vȈT�yϗd�][�c�v\�A�C�K�&��yM0΢h��D�Z����K���JIzNP�RHg�p,�S|�01Z��TzoR���Qw�QI���3�7�ň�y�����^₺�".?��y�"(%)�3�Ă��+� ���f���ؒ�Ȇ�}T�Q�zT%�L(������_�߭�g�I��J���}<|8�r�	���l�jvƦ�^��O�=�8Q��Ԯ5"��t�y:�^����=�f8^H���r��e���5Snp�9͗`�.J�V��۪��JP	���Rk�=�yF	�s�ٱ�r��� CK����8��0n����`ф��)+�NV��qЯͫ�`qQ�����/�4��7�@��B>�*>��!U/Oa����l�DHy����D,<�g'4���9'�B�c�s�����A��|����J?���k���-��!J�lU�L�,��ʡF&�e	a���6u�]�h�����ڬ2kP5��RFg�R���D��_��8a]o�菝���V�/�#��u������$ ��5lf1gBo��\�Ǒ�a��]��N�_��Y�,ҚJ}�dB�4�!�g/^�^���v�׫q��u�(��+eSE���3
D�nC�о�e�y9c�l�=u�
�yc��C�;��j���T9]��A M��t�І��4��YŚi�kR*�R���(�w�ɳ�	 ��E�B������>U��U�Q� �<T� ��~uOQ@}S*�6�Q{���K�o2���C��Ip��>&���ς�E31[�2��
�So�;f�Tb�Â&��/��3�$N-�����	(�v��Si�;*l��,��Weɣ�ˈr�Q���GPk�X�r�̇���������$�P�OZS����?�<���o��7�@�m�ik]���<���+��l�2�a����%D�h�z,{磲�l|ť�b{���%�g���A�D:y���tcg|���E܊�>�:x�/���A�M`����6�/���<����,6����)�5)�sS��`�F�.~��h��g�KC/��	ze����x�H!��~���v��J�,���~w��hj��1�r��?~##�{�)��ňg����T0F�7b� �9��]m�`��o��V�����i��<�!�9�)�=�2�e!�����"\��������d����]�
��f�}�V)L�?������?d��6ף^.|�
d��g!�3��>"�`u[3@����\QAa5B|J!���7��	� B�]�x���	@9��J���(q4zd¦e�?ؠȎ������~u��9z:E���_CaIʨ����ܨ�r�"��wT��Y3BƼQWk=���6ݗr��"�jY�y3W����ǃ�,���?�/��7W牄Y��.x�����w��5͖T�>p�e�}��鋺_`��N��:^d]-��ɅP�P�&����*ڻ��$;c� �a����*��YoAJJ/��J��mJw����{�����<�qQ��St���<}�q!����s2���"��X
��mR�|�}݀=<_�iSbHw�e��(% �K��!����O���Y_��'T��ܕc#�ſ$�b����((w q��EH���i7.��ݗ��ܔ޻�����	9��ӹ�}�tdg��H^I�����*��-�-��uӤ~�!��]dbm<�����0�BF,a��7�"�}����H]�A�I��k�o���W/N���2�O�CF��O�1\?�&e=n-�����X�Lo���r('�����{�/p�c*�0��,k�|50<�`��j�:�I�5jȹ�_>��L�'U�٩w��Ȼ��WI�!�����1nJss˕o�g.�p�(��0X�����l6�YDJ��$Vu$VO�)�R�β��X�^f�P+k9��9Ý&*�Zc\5�;�2f3-�+�Cqh��O6���+��/������}Q�`y�dx�c�7J	=��$mv��n�v׬^]����|�$���e%DT�<}W&g6B���Ʀ��u�z=���v���ɗ^�K���s&��0��& �\�b����� �u��}�R��(�_���7cLQSFcL��>J2{ۖ������]����c\��z̏��n�����,8q�^����f:�K=8L0Z�\�q3�a"���q	��~��!���&V Fs� ,�����#0�������-ֽ�*aŸ;���)e�� �9����@������GR���7��Q���!���aD���6�3���[�B��b	���L��2���]׫��T��e�XbY���ӭ�^/"{9��Yj�In(�A�'��''"�\�On��t�Wt��`Υ:D��@�1�άR�����%�?��f\^k!�a@~0�� ��%{WZP�_U�Q�����l9���7�_��z��O�ww8�����$R��ٵ���|uys���2�4���Ψ]%>���4�S�.:ɍ��jQ�6��=���:ü����w�k�՜�Rq��D�T#EK�W��h��{Q�~���.�m�s�啀�^������/&λ5��K3���s�c{�A����ۢ�##cv�_�pK�.4z���i%�Ru�c82�V}q`؋�UK���D﷥�ب!q�!/3�d̆5]8H�|�C�ٓ�}SR(a���%��TD;x�!	P6�D�d��c@���Ob<S�hpL0���]��'�o���	y�xӇ���������l z�����^�/o9T�
�!6�X�pؒބSQ�@����F>	��=N�ֶ46��8�q����˫���AIHF�VupR2�|�2s-�T�`��]�'&-�&�o�9�a����ת��%R��O��_S��@�	���]����y���ӓ;�3�bl����;"����8�5��<���3g7������>�r��7Y/��u�W7W0Kɵ��:1P9F#�ٸ*Gl�}��)B�Wꊸl�g*�0�~������s���K��v
�U�/2 ���Cy�S`�ILI�(a�?MoA���A�a���)��<E[��+'l��� ]t+S�Ks���D)�*�v0<r�@���2s��x���H哛�[���D����%�_�Q �c/���W�82ܠq��ӿxI��Tk�K6P�'l�X�ͳ�_��|	��oc�g��H��T<bP4�6�^c�����L�.J���W�݆Yt?c����=�9V	�<c־v	W�|4�i_l�C>�]��?^�8Oi�Ik���J��O��q'S�n����Rҝvs��� �J�@8��(7�����P1.{mJ�
���/=���)S =�*���#Ii� ��E��y��a�����*z!�_���㟃Bf��Ώ,>��\v��O����<���I%4~��+��mp����ZA�8�[�eVtg
BRn$g��E=���>�ăEzFy^ �{���uV��[3���@=͚[F\jH�L�\��	�v�%bQmL<7�U'�PZL���E�e��Hp� 6��S�+"5��������C�k8�h��Jt��}���:}����B[��J(�
ӎ�!OA���I��J��T�'?�j��s��}g��Z�T�*Q�8��E:�WC���_����JN�����Z<�'��z�ѐI�跄�!Kr�<)]�
�*T��bc�N���	�T^��!�B~�+��L�ž���7�2aƤ;ↅc̘�
��_n���t����,�g�V�t_1��$�
H��E_�`��$��{;�	굩Z��X2�X���h��H�hO��t`��]��5�}�Ș��zx_��%��;I��!g�NAn����� hS`��ճm·�JV%�
�Դu�\�
����|ZA��.����sC��I�H���5�Vy{@�8}t��4��@)�N�iY���,#oW����P���l����E����>Q�փ���G�S���7�g�#XI�9�`���������d�jy���;�t�븕o��	�W�ԇJ�ϴ�r+��t����nL�^2ZG�OZ �cP$������]��'��e�E�1��	�������5����43{ZC����p�ar�ƍ:QmŜ����
v����NP�U����"���]�wJ�=,��)_�e�cUL��8�u��er+�)I�z�Ll��hYQe����
��#{M(����e����"�i��C-�|�w�y5�a��J�� ��!Jķ�����i��엌^CȈ�d��o���z�nq:�4�T����\��v�-彶ܻ�^g�O!4��j������ 5�Z3B�1Ra���86@{?j�Z����nbq�Mk����ϫ�z�"����>m�/��pud:?��-5t�:��k½�E	��؟��ב��!X��]�+�]A�go�W���2jq?�C�S�d�|Jڛ�$����ӈl�+��2v�z9�u�I��~f��+�#ۛoƽ2q�o/����/t��jI��-�?���^C�� e(�o�S�@�JM�y&ևO�I���qL#�K��cuPU#O�)����x�j�	On';����CH�0?d���H�E!����?\؋���U/sc�@ub.�;�,�R=��n�XlxV64EB    fa00    2460��� �ę����\�x��$�
֚�8��/IĒz���fz]�[���W_����,��Ο��*}�SCԸ�ܦ��c��
��)&՞ha�=ܤ�?T �Q���cƷs�$�DzF*���[�3X�f�:ɚu���!������%J���ۧ��Md����4UZ�����p�˥�b����xx�j@f('�Q5{!�fGCT�N�FZ!��7�]E��P�C�? ���g�
( 4m��[ZϷ�_$��r�$�DƠ���ws�*�9���W��K���!��+;��q���p�%x�zRS{b;/wptx[;m��v��Arw��)�߰�����d��~Ӿ����*�:3l�R��ʚ�B�p���;K��]ĝ�e=���}�̸*�Ń��6O�7Y���,DX��l�Ti�����v-�vt�5~W|~�Y��TwDf��e�4��A7#�,@|Ш`�t��6D�u<�΀�O'Z��\��Wu>�-T�nD����`$:�ۋ�N��J
?� u�'"3��m��i��A�O�<�,���z(�	<Ic��o��֋�K�i &{�#e"V����z=u�� ?��e���ZJ��7�+=�f#���y�[+ޫ�퓔xr�Ŭ_(L��MK=�l�p�>�ٲ�"#H��@eT�$�)��`��W����U��0m3zK��}��Vg�R�O��e�'	��U=��hY����5�Z�{VPPE
��8��+1Xq&��R[�CU��Q  � ^���hi���I��>�i�Fqcaq��1��5h��(�F��Og�ttC���I��ZMo7~��J+̢p�[9�k�0��\:C���qnE|@� Q�-��M����|������i�������]3��|20���K5��Oni[T~eN�7}�S��H��mVf�7 /jM��X2�gp2 ҳ�(���'�[���`�bW�F2Z �σ���{�|
�V��9�U�Ǧ˰N3�8�T��7EJ�I;�&T��++}������Q�1ox��D��Ǟ_���8S���>lxݐ���_�̥&��U�\(^���4�8���lgZm0�f:b��v�2�8���%���ZMS�2����A�#�(���>W�ы���z�+j�y�#A˪^�f�hG�	ja�0����n?dac��� �\ӵ�ux�=a<u��:f:�v�LF�:�� s��c�ڏ��*u�l�N
�H4�*Q��ݒX3{X�v���b5ÑDV��������g�
rV��>&��E��Xk�� ��m��6���/�*�T���Ei8������CAa�$ft@�M���ӄۡ9a���YS^B)�U�z��~������ <�}���-.QfS21�5�̌	����	�(h�}1�&�$���]1y�	��jT>B��|ƒ�4�Zi�˸t}2�R1|�4��f�X����ռ_��\�|P�_��+�v��x�A�zC;�L�e�ЎF.��_�#eV����Z.ȥ�9��V�߈}�v�L����,�� H�,q:��T���퇰�q�����I�MK��>�F!����b�&��,�[���Y�H^?[���SR�$2�2ee�1��\��&��SRB�������"U0;�� d�g������/@��8���s��bENX�S��۩A`�#�z�	�P�G�8MD��k)���8F�,�q�l�	�_��	�ߥn����|��<C|�BW�v�^��΋�����
yK=x�zk�*�X�m�L���mx�!��*�øb���|md��I����NYz��@�Uy������'�G���4}��O�0�X:����$ߘW����ibn�R!a�8˺�L���e���=����̓�=O/���������>��yK��L$n��[�\�w�z�~n]ruI�B��WC{���:����?�HH=f�E 2�Z��5���o������aH�����z#9�}"�G�ά���4��
�l+�X��H/���ͷyҀ$����w[ 5t-y�<�N1�:{�d���
�U���)d�q����x_4K��˨FX&S�񤝮��b�OY��0�4hWF
$�y�����6�V�n-���(&��?+�n��*�g�9p¨	NN����\�g�C��3�д7]�{?�Ј���u����cj-�Ǆ��K�{zkTUD���巂��}6���}R`v���|Zq��X]���(S�x����q�$�f�~��#/���Y���(��P��%9��7�(�ɦ��j�C�D����DgΜ�5'4�w���&7"Sk1��0�??���"(���q����6p!dRߥ_9���K�L2�̝����ۻeR�{W^�=`oe�4��s�b��Yڡ��4p�4�l��_���ԫk������k�nဏvY�
�h0z�7Q��驧����˜F'�B���gB5��2|@Ya���8�4�����_�i�M���!N,�b����$�U�[2�֜�X9�k�"�y�تJ��8��П1c��?�@};��/_]���ﳁ���6�P��_9��m1����7a�gV̰��{���0��I����+��f�l0���:��+u X�GHɒ�磜�L��؍b'��ǋ��8.��`�	���X�#���9n�~/=X7�7c���qDG,ھ��D��Z���#r���^Y.����@1�7�z�
-rK �Y�����u.���~��x�K̞�	6@CQ_���2�h@��� �[�$�H��H- �Ł�kҌ{������wDeÖ�~����ĭ W�0�o����H�kL'�KNJ�fO�.r�B#��YW�p����O��rk��%���l�4��դC����Ы��\�rL���%�%�/�mA�i�^㰪�p&ݚ<|�0"��<ȫ����b�ed'ە?��]�ߍ����F�胡_!�늵?9�m�}_��	!�:#���(-"�k�iSM4��_����'oi���.�S�9q �:�s9�.�� ���Ē~]���-[r-ʂ%�O�W�����
��>͑}ܕ$e�/WY��>P�w�J꼲�b�ʪ������R��Y;'v�j���~N�>�9�C�]I?���n���4vm]o�� �N�/H5�8aZr�N]N����4���h��2*4~f��6nz��R,��QG|#�w�J]�4x'���~��܄5�����{ƀ�����}L��� u�J�R��-���^l�O`51��)Eg�_�;���6V�
x%c���\^1�z�G4��K��_6O��2z7�� v�1�9���gyi�^�=�'FF��߳cM��y���G �S01�E�\O�����rq������o%�����Ӣ����_�De�O�	.����xAz1!8,�j �'��>�'?�<�;e8����������S��J}�����eY�ʝ=�,ܟj�q��S�3E|�p����v5"�fb�.��W/��UN7���`*�w}]�B��mA������NXE��_���G&n�"_���\ɀ|�{Њ4=v��EP�� �m�����'<��^��@l8<wAk��lC8���ЍI�;�g#vS^�7�7�B"~�c=��̳�0d6��O��$Q?���fե��E�UZ7�h%N��9�����p�KnS�6�d׳.c.G��	���#Ua<(�l !�dOƎs#"���s+⠹|������7E<�,�?;Bu�t�f��q�'r�Z�k����|,n�9�kW{+��>�i��֢���__<O�c��bɡ[�B3Ņ;GP�c71Po0�%a��Ae_��v�: ��X����;�f�Om�g%�뫶����9����@�P!�Ɏ �6{�ې~^��}>���E�[��dK��(��]�.��g��ϗ��g���ޫ��qh�t�^N }=��S �3T�_=6M0�)�4fB�'ࣥy�l��.�<��6tB(��>�#M�ԍ���:��_<���Z}��
�Li��u�����M��(x�%��ykV�I����Q������]֕˦�x��+ȣ=3YQ:�cuA�t��i# n�ۙ��Y7���k�7FcYԦYRls��2��ګ�q2��QE�<X�q�.����d�s�c0�v�dO��65��<�du	�!���X���#�w:C�î`��h	����;B�[ t������61�	��{L�����J����@V�aS�m�-?^��q������E0I�uK�"�"��kRa�ң�R��j�n3�ހ	�v���:��Pc�n5�
m�uɨS8��z�;�}���?[��c_$2<B���3�ȗ�)�3~��l��.���ڛN��5'K�k�����-��O���]��|�qK�<�t��\�!B):G9� u������v=�?DXZtC�S��6��L)��$��o���2�{X�?x%
����*���"�9���k7k��3�}���!���g���p���E��1����(���u�%BPp5�1�dY_�M���Ig��eF�rԘ/w��|�|�T�Մɳ�;h�Is��n�ϧ|�~5aUd;�{®r�z��O�L��p�F��qu���J��{q�)��d��*ڞ����t�N�1,����)Q �W��B���vڜ����/���OExT.���m8�5	�|�{��h	;��P�e%`^�l
q��X{��y�ČgkK�XUC�S��:w}u�N�bN�]/�G5�!72~V�����ESa�PQ�Sv�j�̈��(׸�3R>�I @:z� I�V���XF�7d��$~�%K�>;~�h'�/S��~���J��xC�;f�%�Z} ��{��*)��zJW)Q�/����g��K�b/1p@!�I-�6�D��r�V�y&�*�4�f����� �+�8�e��t����(J�\!�����BW`/�#k�gh�4����7�V��̀7-��PH�g,s����ӓ��%5�Bs�rp�)�,+�AMX���+�&U2.�Ek�l��`�I_�B36|	�r�$G�� @�|�*c�f�>��bK��nty��؂{�9�8[����}���<jHN	W�����9�:m=�����~F�0A���	���bE�Qe�����72W�cX�q��@�� �ާw`�,�\����e_)e��$~Μ:�� mZ���!t��<����.%z�@����K�Io\C��]R��(܌���*j�:�[ej��ˈqt��5̞��U���+�y�L�.ꧣ`���ۥ�m�u�r4�[����_�ر����&�l��T���r�����[��a�N���=%�@�R������o�{v�e����f��F<�h��!X��͍����|�C�)�U�9J��>ci^(��їgXr�mr�¸W�uB�żl��Ζ�j��"@ͭ{u=-�`q���ty76�`�����D�,��J��	K���ZN�1�a�%G��d���xM(��L٨nbߦ���d�$P�?���5�Pfz[�Z�u@<yN�f�H��7^�T�CC��{2S�x�D�����C��cr�Aƞª���6�Ľ�u�r���t�o�޺	l#'�ߦ�;Ӌ�����O�[a�h�KpjR��G�C�\��]?a�O�>��2ԃ�1�f���WK3�t;w@H99�9�yjLe������{k��X�m�g3���=��x�qҘ�E�<�y}��������vW3wO{��ŉ��G�0���H�-�fT�3��'�~�L�Y,_�o!�E��VxsF��&���*e^���<�0�b��y(��Z�O8����g�.	�M�Q�<6\8��\X]���������>�gI��N5�>���*�Q��0���;�X����1?)����4�L�Wp�?�]�г�Od�G\�\��7���؉y�`��l�}���p��'����z�ͨ�v~}cd 0�r�t2��dh=� oܷ_��{nNEQ��t�<q���	�Ϣ�ǙX[4QF�_��%��Q/������с�uc�vO�D7bHY	ꆏG�j�ϡ�% �e1�e��9�Z��,=4M�
�3m�v�29y|���_s�����	lS����(B��m��KC�1k}���8m�X�ܽ�]ዥ2D5H�<U/�״�k���>0��<!oLۇ �p��,�l�V7o	���o���rF��ۦrܑi����'">�B�P���sc�{���cc���Q�a2W/��R��Ġ+�2M���$����z�}�^�-a!GN�������^����1Wވ�f��-��)�r:�����"4u��4���婸�dJ�`eƢ��P��l>b�V��$wL��[W�b��
�ORDΦ٤���p�Ju0PrCz)L�0�\78(�@�9PG��T��Q�G��K���Z������+��ߥ��>N�X�H?`,@��"Ɛ�-��*��$�j���-�F�\ty��S��0��.���������o%��ط�+�b,�ɴ 9��N����K�&,��6�ޙHS3V����P�����!���\������ͳ�-��>���������"q1���!9SvC)��l�W���O�  ��'��*ĉ&I����ZҤg�M��C�/SE��Ē8�;p�kL�/��s�	\Mw������g�u�~���yL�΅�������}c��'qabr�&�(��K\�42����s�㻦o��Gy�.�����z��'��{��2Xַ�;z�+��5��s��ۿ���-*��5�U�WN�ǎt������T�Or���^�k�z�L(�p����݃T�g�O|�����J@v�ɫuA~��x�e4kaK˔���ٯF����1��̪�P�T�q�"�B�}Z�RE���.ҵ����d��z�5��=�߅�X7I"��~�ܪy#��Rȯ`%н�*	���"$3��A�g�g|��	{pE��ݪL[TK�.�m�s2"� ˩�b@#�g3ʈ3D#]��+	�ɰ���=m)�)h�P�e5��h}t6W>��6��qM�)��D��5��Nf�Ɵ�'65rv�44�����pUs���F�7_GGpUÛ��zZ�\u�_�l)I��d?,e��5�\I
�»�R�q2h�g&˛�se�Q7On&
7&�W��dr%�V�|M�wa���N�儻m�0�v8	�;�۽A��	��e�,��Yj�"�V\�6WJnqȕH���l��M�� !�,�o�$�x[dN�1іȩ�U��K?P��:4������n�?d�/�
Q\ʩݜ���H{�w��!@l��vm\D�j��\�v��t$5�2mT��E�cR��0;S]FD���S0_�m+i?)󙿟Kd`����m+_v���E��Z;���&�)}ֺ�%��v_A��.�_�N��������	�t�)��m��1�F#d`iH5�xrYg��4���'��B�{��We�,Eە�ۘQ�B����xqqߩ�C��'0�U.���s^�)c��Ӛ�W=d|A�nv�eUK��\n�=�����.����^D����N��7rX$i5՟#d�A���E�H��Ǒܳ��/�ѽm2���b�rDܟ�le�=� �sH��M��0.q�g1��yU{���N�N���Oe�����ҕT,���%V!묳84V�'��i�b�Ν�1���jo�T�P��N�٦�"�J�+L����(�DM��&^m��h��ы�HN���a��WN�������M�.>�������	�G젗[�4��{]��PmfUߎ:%1p�'Ft���:ɠ�ROa�K�m���?�ܥΕ�ش�g��ص��[�_.]��K���P�Hԃ<~���v��'c⯟)�)B*�� �I�x2��(B����\T��*g�q���Fٿ�,5ޣ#��������f�q(dX--�� �{ȣ(�i�Z��*���5=��#$��n��R�{qɃ=Xs��YvB�YaOO
�䡍�8�J���R����W��V^�/��}���j�()�t�*��>
G4��V
�S�K5��98�����H�l��mO�(n���G:"�����f�̓�$������a���S��z�D:�:og��d�0�`���=�bՈvg�ɢ�ځ���w�F���=5|qn2ӈ��Ive��,�z�kd�;m�g�E�F8�u��ʏ�i�b� >Ǔ�0�抔>�(%���P�Ve��H�ܷ�a�Ӳ���(��(�<h�i��uС\j�,v�'
v�(���5B�T�%��&�u6}G16n�m�U�왉<����TlPC�=~���b&�=OZ���� @�X��y�f�#�9��׎;��C:���9?S�C�b��x�Q�̙υ��@������3$:��k�q�d"tq5r��_�,5D��h��d_o�Η��2e��v�m��7d�Ozr򈔮��1���[���!�XtqN��
`�Zۛ]�SeVjX̽��He��R�ʁ����m:,����;�>�Ȕ�^�e�dA�Ԯ���_Z�
�&�����Sp�je�.|��RGl*1r9��򠗬v	��A�|R{L.�����9ߒ��#^�5J
?�%�ew�I)r6H�nƑO����|��S8�U#��iox��iױ���ٔ�Wb�!���j���`^W�^w;�*O�К%Z���#�9��A7ce}��Z��<c�����C�抩����&���]� ܙ���}���n��=ɹ^�35H,[tf����lm�+��6��THUu���F��xL�7�h�W�"��xF�ÚvDF��ܟ�xjظX`�5c�@�'X$)=���Yd���&�g�fa:뺶C�3�pc����a�X�� �bJD���;��Y3L�Ӝ!�j̴�U2��#�qꕦM���O_k��6ў�I����^\�=����9BFh,v8����j���{̂ݸ�H��S�Dad��w�p���g3sdi��e:.���}�O�Ō7J��՜�I0w w��gJa�a� �w�&��y�[QӘa�2��t����K�P�}�"!%�C���~��9)|ߨ�AN��rB����kӉ��H>��W+�e��Ңc��]����%���-�'�S�4P�
۩�7!���O��=���6�+�+$`U�A��Qȃ��#�X��Z�
�-:�4��"1�'K�!�Ȋ���c�z�u>��d%6�?��6!XlxV64EB    fa00    2230!��������M���-C`u/�Y��m�+m������gH��n�[鮺IcdF�y�I\y���2�w�l6������������K��u�+�%ێ�k��P��_od{�C9M��θTE=��.�3��\e\���w\,���_g�}8�1Გ������!���vfY $��3}>�ke���,+$d��r쯳�.�����2�,2,t�h�}�D��r�ߓMYTaQ����]}
R��`j~���܍?���6��<�涜�эn�&��`;u���Q%-+�'�=b��X,:�Ig4g�ƅx��oUU����uZ�4�B�K�ݟ�>��)O_[�N1"|ҟhaaN-�VT�DG�ω�In�rDȞ��T�8��'23���C`�x��H+�����?1�h���j�e,���74Pu�����G���	~���DU�øwV��kj��%ϖ���k�S��I (����ڲ��"���zr�]4�6?F5���?��kkF9��fKP�!���WY=��\�c��`��S�w7��_H0��k�>�����q��1n�	��G�AaF�`��e��&�]D áE�ƕ@�2O'9�Ө���Ku�O��K��I�&�t��
��hY%�]��^b������	���D��%:1�E�Cޫ��?�5��uY��Nh��n��E�Z���U�aHW���k����{Y���.-��3���ઋi�)o&aeM}PZh;���h��,�# ��rx� �8�FY���(���<����g�V`��	
��ë��1ғR�Y��A{XO,��'�V�\M�x��D��h�k�Qk�L2�
YV����;~t�����=jv�#u*�|&�;a9����P0����E<��}WƮ��j�4Є�SW-����mݛ�69 l ު�O�[��Rt��<R��&_b�<�� v�Ǌ�����Q�T���Sq�q`Q����+67�&���HGc��H.J0��#�Jfvʬ=�	�y��(U��6Eޠ�&enV.����{�P�o���&r���'�"�}Mӏ�Kg�#>���vv'��_�P��}��f��E�͌�5/��B���ju�+�Q�i�i{@�~����u\�Φ�r�s�c����.��N�Έ�aN����`7���@��Љ.�{����\#�,����U�BK��u�����{r���+N[�f՗����#�vh���" d�V]A��ߒ�>8�V���I�N�¬�{�I�4@�i��t�ſ�j���z	��!�1a3�|����A|�Z2�d���V���4˔���
sTl!(jy��]�|,���ݧBxj,�'�gK_]|[���d�ƙ����b3���&}z�쁬�֨�[�&qg![�63�>�c��̄z�5��Rg�rFmF���Z)$���v����5�h�<��K�`S�r���Z������=G����TnG�^��
�z[����^%��9@���Ϳ|�f�8�]F�
���x����\�k��Pu��)����.�� �2�@��Է��A'/���N	u��K����:�o�����D,%��QJ�z�'�\�Y���a-�R���,w��_3C헅V}�ſˁb�
A=R�+�T�,
=�F�3���sԢLc�_q���j�CN"'��3O�K$����Y4�+1�By5�g��	�����0K���d�
�\H�o)R�Y�}�������#!���D-��6O$�1���j�t�pq'�]���i�����W�34�J�짍Pd�k��g��d$c�Q�k��������EO�^�jK�5} ���``W�b�")��XVUj��1�^�Ԡsc��-f�z®�Ç�ſ����}x#V��Zr��_���۠T��= M�a:�B�
���ݧ��ཾ �g�:+���^A���R�s(���Ó���Zw��1�t���x��G�)��:B(�߀���a����R町���9}ơl�(䑚?��5��W&P���m ������P�EiV��g)ڴӻ���(%�RNY '7X��B�TI�R���Z��r��i>�B�>��\[���*
�y��|�*a�cv��Mn�����2���ŧ���Vk��Ϲ�����HB�3�S���"CI�	�%����ķ`�&�^
�R��BӱN9��
Y��繃��x� ڿ��d(�E9�aR7Xz2]괆�L��}t"$14�S��	��;,�7cg+�)vn,*��f�+$�Yg�t�m�X�L�@Aa@1r$��:` �}@��d&�H�#Hk�����3�7��PC>+phe?�x�n�4?|�i��kN"��Rs�v��:�9��^�48A��Mk�:BB�./�0K�$B��N��8Zb&Ǩ��Cw-��KF�u&�!
 l�z~������_���ͣ�g��3��<��%Q͎c�F��z�T۞svΎJn�H&�t3Z�6�����fSc�aA����0�+f�e����gښT�Ht�����T:��D��T6t�Ga�h6]�sR�_�4�����#W�zu�0�������6
@,�g���Wp-��5��sh�,h�D$d��"�uY�g��.�^Ocd�8s���@�1���v��q�7��е�FmW�8��P#$���"�YD��Oߞm ������;k���/� @w�����c����e�X�7L8k���3��S���]����h��C�Ý���[�m��-Rg�1�'b���"ۜ��Ξ0j�V�T�w��甫��ê�B��a��Ht��T��6S:s��e�"�z��	.��H�ϞvR�e�P.C#(1"��%��hZeeo&KԸ�����������k*gkh�#�}�Z �X5�у[�ʟ���m݆��㊤9�1�HH�9MfAt	~unmN�G�,�I�y\�<�8�5&�~\V��M�8�It:p�fg��|�뇞�e��ͥQ�$;�&"�7L��PHm�	;�b���`� �F�*"	����/�dmm��t?١uT���A�(�Bb��T���w��{9��1�u�#�<���IJ�&��C,_Y�S�� �ёT���{��U;w]ψ�.C&?fQ���Z���P��t�B��w���Os�,�0@�:p�?�S����[E��#�(=�����6�q��p2�fҍދ�s8���a��֮
�^_mu��!�A��z�*_
�|�C~A���
���(��q%]�Jqv���b��thT'��'�0y�/��2i|��^PC/U��ݏ�.��2ee����-�1�ۇ/6�ǣ�s��W� -���,Jq~R��q�ͫ\����lw�Y^%Q���I���[J<�NԲT��]����TH lQ�ѽ�fX���� WA�3����O1��d4��l5���`<
"��A�uG�\@�X�7yn���Pߘ��'��Ø'�%U]>� 9��J�|t�i�<���C=�Y*�a�Z��J7�����)���@�Y��z��sӫ!�ۯ�0�Q�Rj7�H�x>w��̊�{�����B�Nev�Ògzؗp4w��}��_V�#�bp�:/G�5�CwC�p	m��j;*ځQ���x�"龚�6��3:��b���wX�~��MK���CB�9�G�X}9�W�ݤ�	�������I��F̬"e���
\L,�^-��M�N�aŻ��E��[@ic|z3Rl������r2;{����)^i��v�� 1Ǔ� 2�Ǩ�,4����D�?��\��븊���=a�w��܌}�x�&��7�җ�r���W�WlH��Y� ���a�E�ZUVv -����:�$Y)7���fߘR�cI���<ڏ;���LĮ�YJ�����4͊5���'Up6�p���໒��w�"�Kt5�kݲB��f�2����sA�/pZ�B��g�,%�����k)��rH�kS���S{qT��~;5�GI�Ӹ�}�T�q������
P�n��I�1�=�}�ǁ�6�hi�'����hK�`<y�Y,�ճ;��Md֤��Ϋ���
�o.tJ�`��?B�X�A�HI�ݗ����eS��	6!TO&P���>�����U�������!����������8��UR��*cM����/��u�Æi��s&�w��F�^��)�q
*X�I
��x���	u��������D��l���8��o�!,�U�9�=���.yA���߿�n����"�:���f7dՃ��JO٬�@��y�Dq-���E��� r�7�(�D��A���a���h@l��5�;.a����'����=�L�9��5 �4c�li��U<����Q��\�K�
j�ȧ�5k�����:��B����EFh��s�<|;��ʨ0�md7wU�¤bL�ŜS�6��z[s��f'�ۘ�]��]h�/b4��<�uQ֎��;��^|	f�Kՠ�I,�g�Y��e�T/2�&�3RZ�hc���#��ִQT�$'z����z��c���m����E�1�i����%����=h�O�<�[�����'�����95�H�?h]��rv;�,N�hWi�_��i���m�$�d�K���e/�}�_
��F�/<'t��p������|�L쳆�B�1/IyVb���/bf�!:�0km��7�R1JT���h�ĠeE�$J�4�S��WM�Ct~���&h^{ǲN�o`����#*���5<m��� S ���I^���{;v��#�*x#�=��l����-��@�rZ5ʈ�+������Ro����z���:��$I.���Ժ}$��j����
=_~e�Vr=� ɑv�����3�;l��Z䖗�3��7
|��������ڗ�Ա'��H����o���z�P���e�"��-.bUw|�u���crf\lo�,g��v�U��g���71	�z2�r�-d�)ά��ch�^�����8�ZY������ʯ�Z���DO���vy��5h"��<��������6֠����1�rE�,�r�G9�y��0;��w�,��f��o	�r�r5���F�	�t����"A1���[	��m����?�L-���>(C/4��s���H,:��{%�}��(UW�!�P�/|��ʞ�v/���,'s�k\��|u�B׶"B�=�����k��!�?
x��o>s�Ar�IDn�L0?��J��[19�|�c�G�"vS�}ϋl<�*UW]�L��8�ۧ��{�"f���敡�j��� ����RԎj�F�z��*�$N��cL|d:�Y��}y p�F��ң֊�V���k����v�ZhF�S�86�_�Zܪ�L����~�8���crQ��;] �-������S~bUD���i5
����5V�k�`o3�u���+Q0����|�Ub���<��#���=�8��a	О�И#�2m�ü�m��<D��R�Կu���#��h�;�(�0ʐ(Z��>�D�T^�10O��-�e�BP�V֖��E&��!|\E>,��b^Ǽ���!Sgфge�Fr[<(D�JW��њW�{gM��$y���F�3��u�e�HB�Ϟ�r��7��H��c��0��k�fs�f 8�����'���l��o��i$$S� ���M�T�Bыd�QP�Ł������H����,lR2�+ *���d5\*���X�Ǫ[hev��7��<P��j�=-�sT�l�D'1p�ʬ$BRW��/r
`κ��{!��=-F�s��? @,ͤ���!�@�\P3;�{F S P�I�u�gVޙP�uw.�DO#Q2-^I�n*�c�������s�P�qro �&3u p��x:�?�l�c�ŭp�
\ST�C�YW��3Y3UJVde3w�h� #�m��Ez(9�u�Ω���A<D��8"�t {;w�^k���w^��A���1�N���.$=V�t�T9֢�!���UfD	q1�X*��"�*��i�������� �����z|��:B9�W��
]�",�R	����i��')�N����upQJO�Sd	�����(Q/w#�R�n����7��f�I�!���j� [��%���MG�*S�3�iI��!�����'�s��9pU�EkU�;��H���T� ��� B�!�p� <�U����q�mZ���yŢ���ժ�wp�5�>����� �C|{��o�>�(/T�7Q�7Q��V
̥�`B���f:EMb���@�`#���j�8�]aY�R���u��s�9��?�yG�:$��ek��b��Q����tZ���!���g��@�:���} �4�],(!�+�v%B��rf�C3���tJ����H�廧W�����i�jI#��sм�0j�G^���}�Z@�Ү����E�<��R�1�0��^�����^��_�|��+�a���!����W�9�E���XFn�����!����Q�ڜxS�/�f�h��I�D�s�rds��t�?�x�� HS�,cռV�o8��EO`�x�m6����x{B�x��\Řy׶��J��i��m,b��d�UW�a!��s�y�~��I�I�
�P���Ep;�x0�C}ۈp��_�?#�?����A*K��.��T��a���ݴ뒥E���y�C�cn���(x0�{W�����c%X�s�nUט�_�x�,)u]�-o�2�ϓL�GQr��,�0jdN1�6�q�;ED���pP�+�E�������ݘA<Y�O���+�=1�����s�H��o��L��,��DW٘���T����P����c#�!o�Di���݄��U����v6�է�z�yS�ᗪ/;~|p?�n��P�=����j�Lsꀪ��v���P��:�{)'ĉ�����K,��~����酰 ��^B&��ԙ��=<��63�K���%�aC)�S)��Y���ŕ	��o�=Y�X2N�
V��u��)O���j�KC\�����#��
?�zO��y���N����q@�e��}ԏ����k�����Ej���.������4k	���`�?t~Uf��1�)��ѭ�P��?d��k��A��K�+�(�GGR���Ėrhr���4��"�N�6eT_�:�4���*֗�-��3�?<@E���]���h�� ��[��`E-)�Z��e���.�ęan���{�>u����I��0����W���DZ�y�D8�y��{ȋCM(����V�׺V ?`��:��3���h�0ƣPX��is�}}Z=Vlo�4�m*�h�����l�����|70��9��KQ�q����)u�\/��0p��Cf�˩��+�E�Jq�
Ҁəһ�k���|E�wz��҃���~&0�Q��T����q�,dC*�ny�
g]�����ɒ����蟥����ܣ�����������;���q�c��ʲ��U��%>��1�;-E�Ɗ���P���$@#<�.��w�3�e�R�S��|}ka]��6���e��`E��CiQ�w�<��<���Roе�y�GG�	�οtKk�Qi���]�)�袸؇`����wou�B�e@=�q����0_�V��7K�#Q�)�5D�����W���98�׾�Mۿo|����/�^��aL�Š&L��dH~Xb�q.b>��7
���t���x��Z�Ŝ�/?�.7��G�[� �:�W���R����9�R"��{�e&�B��5k��#.�x<�@^m�u�@����Q�:��ˡ����7Z��f���WH��!ְ��� щ\�#�}�H����z����,�E*H�/�L-Sh ���q,V�)�2[����.��x���3=��FI'ݑ�Qu�"Hڔ�����	�c��ՠ��0����	��N+Z�����>͗_6���˨�T�'��]t�2�l��a�R�
�6��PF�"Ӧ�#ۼ��/YV�󚜄��a����8��o)�dX��X�=Ze{�ps��:���A��k��
=x}�|�o�����bLی�������m=jRM�!s��2l�2q-��z1�����ٖ)��M;�c������AuP���-y�Uz���&=�Ѣ��i��L�y�ğ��-�&W|�lb;����v������IҎ� Ũ��� ;�������G+���M05��dIdNt����T?��t����/�b�u�E��(I9.Dō�p�7�!`�bI�E��Fn��NJ`.
;I[RB��%V2pNU7��v��.�
�s�)rq�$��ͪ�(����l���ݭ���[�U F��p���M(�6@,��¼p���C���6B�Wj�Ճ3Dn[�Þ!�vf�0���*nl��x �_���^hu�1��g��9({�ֽ��;��K�����^�95�NJ�3Scڱ��ޚ�L��\1 �ܦ�_�*@jZ�6�|�l�w�֧T �B�|a�/㄰ w6��|�����I�h��{|7�/��d@=��I"���M u����i���"��jo&
Lݛ�� "f{!b���ب������]��C Ϯ	����jᇙ7tu�:��A��uh��$	��wPUZ�{A�I��WY�x��dN�A#o�HdL�ͷQ����K'�F샠��b+y�����ўH��õ��ˉ��yS�Y�x�wҴN?S�O��ոCXlxV64EB    fa00    22c0F:������Kۈy���#�?�z� .�;f��\�ܫ�TR��kgݨ�Oٞ���Q5C��]Qá?��Wr��@�'�YՍPM4�4�J|.�8�?��g��ʜ�݊�U�����:An�;I��������K(*�5��旒(���%�P��&!�J�=��ݷ��ڣw��M����B�'a���ن�m���7V��
^A=�$Q"�j��0�Y�ǥדmE�t����XŢ�o����[$d�G����'�BX�������s�o��Z�A�>]�M�%��"�t��OC��u�Ph1�E7�#t%���QId)!?Y�狓g���m������G�rO��d���	k	���wn�Gnp
S�]ӨT�R��+F+"�P�{���m� ��}|���[N6*׶��xߋ,Nn�&��G��MqX��r��j�*z�|����ӝf�k�qi����'�>��F�#5�z�j�%���5,�O���i{��D(��v���V��_I���T�aۓ�� ��@��r��n#B䡢'r�iKs����g�4�����v"QNe�q�ٔ*|�������$(N݌�m���LC��˹.b��:�{c-��o���H�7S̸gͲ��V�C�[v�}��7�T��5�L4���Z:N��l�X����Ė>`e2/��!�1���:�Cr-��H]x7�]���Cx5BN�y��m��Γ �"���O���v̂~���� v�����ڲX��]�?������Mޒ\�����5vͽX�|RNڑ�)�8�s��	-�
��)�?!@��Zp�~d��/3���hлzT}y�ֹ+��w"�
�������~�~����5-4r�e�#�v�u/K��G���t(}��Ӟ7�[����g����~�����
!Q5�]�6Lb�����@��u�/k��z��E�Pbr&]���܈��S��4Ш�򙳺�Q%OW�v�g�,���$p�D���/-ۻ��fG�3�`Rv�j��ԅή̍��&7V�8��H�/�,v��+��/�al(I����=����&�緣w¯�Vj��N�1����!�P*�c��hF)����8�ǧU$X�!�����J82��&)�T��{t�ٖcZ������3BM��fLUc��E^����<3@�p,~�tշ0��ww$�&��p�����nY9�6G�vw<p���f�ⓨlD~�1��mf")�M�Ǳ�T��q��8���>yf�⥗��I��&ű��Z6���Y� �
����!'ܖ�۷�U�hG����Ea+WI�g_����S@���L�I�ؠŤj��[��)50׺_�)]E�����,��7IFE_��^ �ӎ���	����D� �r��:���_I�iu�����,�ioI���?��Q^���َ�R�W�n�R�Fk����G	e3���u�,b�45�����Wg�>���%)�ǜV3�`P~W���wX���>xd�c�Z�8���'R�l�%5"�o�OK�����{IO���<T�4�%���b��U/TI���8�k{�.Vڵ�QʣZB�5�m�`��1a��`�օU4�G����<<׃`�=�� ��Pc�����x �a��
�x��бƵ.��������I��.`�Xfi|]҅��#Qw����n�+�cɓ��~!����*n���X�D�h�[��2P	d����}
���t��k5��3 �BQfC��'ۧ&�JB�JKߠ�p��QbtSA�ͤ wAN)���ݖ���K�[����$U�O���σ�2+b�YqִK�#i�#~xga@zlp��QNt#���&�r�� �Љ]��#���'�Ny�]�#a�V9Y�烌��w��w���;��0��q���hU�x۪�+e+D�NFd��kF��8{fD0�v���L�]YI��� �*�����Gȥ�s��g�,�ڷ��-�ە���P��!h�D�*(A�$6����b\�,��� �į�s��A��=����`fxn�5R�J��?R.77� A�e�V�x�7�Sk�����R�1�uy���U��"ٖ�e�Nta��a��2X�+�I"]3�]�#�V��,@~�Ӓ�ތ�
�咴G
�� Pq����CS���ΊN��ƹ�
㻳�O��c˄�`��v[#�T�:_�q|�q�p����^۵z1���B1J�ׂ��C��ޜ,�
]�L�{*.��%�{c9�H��/�|g +����Y�)��mZ�a�<җv������f�l� ��3�5�L}h��ԾS�!�=�H�.�������p�r}f�w�1@��?k~'�ڃ�NB�ɝt�a���L�mU(�&A�D��_�lF6w����$((U%�~����'�:��ٵNp�Qxp)��-���x �`���{LB���/riNv�Y�X��{n����L�Nw5k��o�6�[�yedlO:��[���Ȩ�^�Ơ��dl��/�sñ]6�L[�8�b�,�N���.>AFE�zA.�_Ŵ��)>��¹].���A�m���:�k,ϕv��!W����Զ��T}��
���z�_%- �z��:E)3�y'Be�h+��C��ն�����(��i�|P�����&( ���e�u4&0#7�Y���3A`����T��9<<M�Na0n%Hq	 3ͬi�g����E>;XK	{�����v�@�v��m>{2���N�{PG=Umu@x�<)��
�-c��a����P�A���4o�]��f&[8��M�.���uK�7z���HMr���-^�7�H��V���P�=Eu�����W����(ܑ�}֥�1�X��*�~��8X���|�2�W�H�:c،�<�ŉ9=�M��6'q��Ή{({�n#�2O�fˉ�_�v���&�#O�%R�?M8J,e��ݿ��Q̬>�SH!xql�=p1��^��WRu�ޫ�Ĺ���D6}0��67Bn1p^�)K��:�2�}zn�odww8<t����%1HR��x�+�����aq퉈�#늊*h��n���6�Ȳ���͟���d�S6��)<�r4_���G10����Y�x_VgŘ�R0��j�d�4g��������}�5X�7Z<!�BM�f?��Z�^��]Ď��4��b�w�ϟJ���f��c���O�;d�B�j�F�&�f�Y�OEK�?ٗT����|g���I�t��6q7� ���S�\C��{H��Oo��y俧k 7�t�,��qn�����j��Uݶ�[�r`��.�p�o�̀`��M�$~�,\:/�aR�@���$��ci��O{R �J���b$�ΰC/S�: �� >TQqv������-WΞm�&IV"Œ�
�PR������_��W+��$7���.@�zp	0��n����-[uK.�C̘B��I�:��&z�D9� �ҫ/�h��G^ �~���ڵR��H��ۼ3��6�����`�\�M���AqUڬ��A�0��� �e��_�;-$��c�8�/w-T�=�Q@�m�y ܡ}�F�&rV��E< ��띎\�����B��I�3���J`��g.�a��sm�$I�1�t�����˶�̵��ԥm'>s'J^:&3�X�q|^��u�xR�u�A�3�9L��ʬ��p8���۬ν�ߥ`>��A�oH�_^�p�L.b�vL+��
`��m�"LB��%sx򕙹ME�yx^B豈^���`���2��ԧ��D��P�7�&��`B囋@�s��lȤ.�D�_>:(Q�d�����C��,TT2�M2��F��lj>��/||�ǅ+����0+�jWi�b�ll��+|ׅ�K�o��G����[W4ѐ����t�n�)�c��u��l��r����	���K?	�eM�R������ �G%���I鬑��j�^�b{R��}A����_4���tǶU"��E�� r�1߀ª�\M�GL͉2a���gO�j���}Z�A��'��y��1�x=���I̓PF��nTl{~w^�pk��úY�Â�a�_j����4Ŗ�L�4�θM�SQnF�m̸���K��W1|� ���HV��ha��qeF��ClUr� �h��ީH{�rn��1����'�����U[">�1�7и�՚ȩ71|�Ҫ=2���� �O�e\��a@R�{��3���~1S�81�����'8٢��sFq<U=g6B�x�^�]������͝7�x�T��7mի�$�qr���c.�t�UñY�{<@�5��Bn%H$Ke�CvP�8c�|�c	*H52����<f�o�����iu�r~�5�4��+������/����"������Bq4fw�����(u�ڛD�vOH@>���ɓ��������cXKP%���S�l%{HEu��O�҉j����м���0���V��~�_2n���E� /)Ɯ��2R�xK1^�T���k{�,�?�6+�b]�j�'�]�ho�zq�.O���>����K<���Z+��׊��f�+
E���\�	̧�7�#���S�E� �{D\4�|��7}v7ip�z
�R����Z��n��d*�눹k�j`ʇ�4/�ݾ{n�^%T��Xyc���UU8{���#k�oU��"t� ����׫1D���"kh��A��]�i`��0y�]�-�'I֟KH^�K��dX	IQ��J��G��	.�N]N�:o��w����;�Po�,U�8�jk�� pE0LL��mH�T�3�����,��[�A4���
&�Fgׅ*����-��F-r�l�2�=n�V��z�܈卩3���iLK\T�h���=	!���0HьqA�TH�2B�t�7��^�C����xA�0C��Q��X� ���oP�	����3&^qTu���4(6s�L�Z6��=�-5��C�M����a�2R��E��a�ο F��eף�H�bi�M-����.G�N(�O�|X���[T�[W{�X��X9Du>ϗP�m[9܃C[�Q�"��k�K}3�~�v���k�-3����h�A96�ҽ�L7zY�f�'x������:5�5pz1E�_&��~�WT$�G����:^�Rr��+�b�A��!Ҙ�!s�H�xd�I,�n����inV����|n�	�E�x/��d�S��Y�]r�x�u�ڥM96���Ӛ?�6����x�Om�D6K p�N��h&>�ɳ��<�>,_wT|:��!.���-$+fʤ�;�׬�g�=��O��M[b7��R�H����hS/�M����y�Õ˻�uDy˂�Wv?"J����!�[��� }��\I�̝[�_'¬�+L������l�;Zp�_��I!�A��{u��L;�����;���6qcȾЫ�_��%��$/Z AG)={�����q�Bq%�ߛ�]�JW:������OA(�p������d��qt�M�:�'��a5鐍�;X���hh��yά���Ei
u2_��C%���:NY���$"��X�@ߴ�sr����{U�0��y���e�0�Kw^��f$P8�����=J��@F�HFx��o�z�x`@�2C�0���V%Q�w�Q��ï�K�e��U��~�E�T�0�#��d��'��Z����Mk+h��'7�>��2B֥�w�Ƈ����Ӈ�чW�ί��\�{?�=N�?�����Qe�����j��ܟ3�V��P��U���O.�[B?XRD#ײ�5d
[^/�D���{������ǐ�:��m|���]�Y�Ւ���`������#���1�r���b��Wm�RE����&#�f� h�2�B�1�R����$��q#�����Vrb�����
y��U��7����27�R�E��1�qu�2��������N�IH�i��8����Pigʾp|�_`ٚV�ð��������)�^B_.b9w��K7�:q.�ڞ\�3��Q.��4�~45����>"���5F)�(}��	��еf\�r��8�+�%�� �:,����o�KsW=����
�j�����`����j�a#de�`�M�po���\��g(�U��3�;k�"n�}�f�N� ����''�ϣ̒m֊���׀��[�Pg��W��3l��,|.6�s�����!5�������š��)�V��D�x��h�P�7�6|��Kj�a���@_O��(\�b��%�������{�#�v�&���������;T���	��u���a���tŬ���rz����o4ͩ'�7x�B�eP!���K��p [�W�H������DԞ]x&��N*=Ɂf:`|�R�i��yşv�>������!����9̐�߳r�@���y�����JB�UJU��@��6��5�7���[!����L�oS9�F��i���
97����{���J:�O���{ӻ�F������~u��N�T"X/��Sv|�V�P��]n~Ƅ(��/���J��T��Qr�H��ib<�h\�h"���;<<��p�X�c����앫���)��U�>悒�CBf�>yɟ�������%fXL�X�Zr��f�.ed�$}q*a�Ȯs ���yߩ��"?�M�ԯ"�k[��J ����d��`y����'sNh2�S���(��m�C��)~]m|;�Ѽ<xTC�?��.]<��֝��ڹ0�b����]�\_���h��X��..��c�1������v����;��]~8��B�	��I�.���XN�	�/���+�+�̈��_J1ш�h�g>�#%� �!R���E�������`�>�$܋���r\��+ �R]�U_z��O�qr��Ф2[���[N�`��C�7��۩����X*b%�_r����I��+c�{K�����,8+Z�.>ob���k
	Yxm7/���ˍ�:4ժ��߃�`͎.�"5 z��U��)�\v��9�-�ٹw��1�����Jb ��ա��x�G)8��B̣�Sl���:pqXBl£Zr�k�Y,��a��J� }I%��8�ש1}�46���ǜ��DaX�����q��������s-�)N.=�ads�Ug����yKfm�3�7�(H]!N���/x��fә�Fg��=;i��2ʙg1�d2v����Wj��2��������딎�c����bb�=鄤gЩ��^�1G� �Z��H�`z�,�,���6���B���ٰ�5F��<��Zx2p愋��Q�ʶx���a�4�,��f<���D�RO�I�}_TZ^��NCW�F�v^���x����f�Q͍�����L{ӶX�)��U�۲=a����Έ�/�d;�}I{I�X������YU���"����j4mo�!`w��N��a���~MԂ�,��i3��@|�
� ��$�둀���0�Y�
w+g?�ɖ�����O)�W���]Z%!2<�BPn����8q{�T��S?`p�$�i�� G���ž_��&�����Y������g�@����|	�8��Jb���ّ��9�ŷK@OE��,2LJ�^pFr>�X�����r�ě���~o�8#
4"-|Z���Z�4�;���1���>ڵ�d��?� U ��ܵ%T�A���N(�6��q8���F����V�H��֥���h^�mz��O�-=�8����ؙ���D�1�����P�6(���.@ Sܹ<�������,9���z��&~�2�d���~�^���7@e掌�S�s&�����>���������{mKhc4	'�:=�j�p�V������j���Ѭ`t��=�&ϻ>#m$8x� �1,�����nNLM�Ý�u���ަs�ԒV���K1'����e
�=}	HyYl��Ms�usj��`��mվ����Ϣm�:H��U�QV���I*��-�r.���66�[�T(/DHu0�1�P��-���spo��bcfA����nsm�
�%F~�R�f5+<ݻ�qͺo�QZ,�����0N�f��ц!���ܬ��@g�z����c���,�D\���Ur7��c�s��l�bɫ[,S�:������I#�MS8��}��H��3S/�v2z�~%ƞ��e+e�NR����6��$C,,raa��Ql���<�҄�s������M3.4��&���`ۙ��ѯ�7�g�-7Q!R􋪷)��jI ��w���l�q�Q�1��nz�/�(M���������S�cIF.jcN��Ll����af���.�&�(�ƌƎFi����&��w������G��ځ D΄ úc�i(���m�n�/��z0U0���cl����9/T�D���i(z��C_ 5�g��S�Dy�UqI��
�]3�Y�A�h��z��5�Nbx�$$q�������Y�h��x՘1T\��rT��ڝ䑙�A]���'2�\��Љr����t.�(k�W6P�ZM�K�Ä
���'���ЩW�@Po/i�t�
)4��a����ft>bj��%�%��R�ַ���<E>��z�V�)�v�f�E���TC|v5�FJ [�B��Ul{G��g*{����rt�i����H3��O䶘�,����p�UN%�o�p0�N"hE�������%z�p�}�S���>�T��a����,;��Z"2dV�+�rՑ�Y"KUq���I��>�\`��x�Ɏ�� ��,���VP�'��|Vm8m:��R��\����@�j$�6\L��LtX��`�����ݏ�f�s��{�=�?�����V��C6��'5��48XlxV64EB    fa00    28b0���_a����:��&�G�YI�3',�?D�aZ���'q#VO
���_	�ڻ��� J�\��3Ao�}O�
��]�4u�[ҁ߰)~��DA��`0ly�{��#�e7���P4諣�I�G��ZܰKX&";�?4K��d���x~!_�d��[p��-��%�Q�R~��{d\�X �YT61� �_ 5�X$���m�%`K��ő��2�ϟԓnD�ϒ,F]TzGa ��o����Е|����U��?�YJ�gֻ]ߐ-'@��N��v(ى����j�J/M�%l�U��'���;@���c���a�	�/���VU�[䋭~�ŋ��;�:.>S	����f���9��ޏ����{g3>ḻ�F��U�Q�WM*�7�w����"���������)���)���˼i���:,1Q؛hM��t�����7U�$ux���B��a/��Ĥ��H�sA͜@�/�f��Ee�L��r|ª%B�a!�Q9������&,�����ihY�j����N��D}4�O\O���2٢	և��Ͽ�Oӛ�	���|�k�����o<z�Ћ4(gC��L�@��oi��5�H�c���;qy��vJ�ڲ3o(�G�?n�R|�������G�@xQ��R�T����绌�o�H��C[�Gz�l��E�5���8���]/
H���J��{�.x;Y���7���
����i_؂G���}al��kU�FD��k� �	_=�|�Z9�R\����M��"	*K>�����"�V���KD99�.2�䮃�?ǉX�U���1���}/$H�Ml��f�Iz���/�`���f�o]����v���=V�gɏG�2����Cek����y����:��9涁�{-?v���_T���qm��}೓L����-����)��Z?�ٹ6R/�O�c��ʽ5�r8��F���T�Y֝��7������7�M#��9��TX�G�I�r�o	l�q�Q#���������� �i���p��/7O�Y������������r�ٸ}0�!?ki��Z�9Ҕe�,T<��y����Ұ��?�,�z�"���S�_Vi�6� �.M��7�9r��?a	��r�ʡ�q��Tޠ�]�R���`H��Tf9�Pa�2�W�0�ʜX���9�ǂ[*��Ә�a��!������*ў^7d�qr/c��I�=���n7�S
Ct��L�g�C���566x�{=S�x"	tQ���l��x)�o%�	v���=>��ޛ�{�˭���Ap!�3��Jψ����)᛽���_v?n#�0t9�"�ڣ!�8��O��&qvf�R2a�vOjI2n(;e �_��V;����5u����PF��=�vʹ�L�DV%�x[X�BQ% ��j�)*}�O<6s>�F�ÈVG��w�1�̒i��ss��q�܀�?+�_S�5��VP�gpS\~s0%m�{zV�or]	Ɣ�T�3MZ�G�^6�m�N����P�D$ރ�u8�6��a�)\�C�n؊&�5�d�o�B�m�����S�@0#�΁T\!EIvt̍2�\N��Gl�*��E7�W��wĘ���"�,.���j�1���
����ɸ�]�J.c��m�u$��H���=)_����<�ݩ6�59�<$���+��MrKqG:`�`�@��l���i�yy���v���U��Cf����0wR
���ȫ�ґӈ_�y[1��BD�\r[�s&�&���67Ն��/��nL�� sO��,��k���o��(,$ֈ��+�<e�fh���L#�
kc$�Q�Ԡ�=������X���4��]z�p(5��3l̣,�l����N��P=��t�u��nv�
��:К�NxX!���T	���g.EHv�/�Z$� �f�:ñ����������!
��>uƻ)>�D�Y9�ܨm{��`M�� e�#tkxjޗ�����<����5g*��*̫s��d$���SV�>�lN(#�,5�2��L��z��Zr>�G�<�U�Y �I!�|�� 3C�Q�Q�(}�
8� 4�WQl~�1ͷɶ�!eu}����3��ꄒ!�v���
��W��1�����&-�8��;g� ���'<ߋ\'������^�,�Q�[ �5�0��t΂�)��)��I��CѮ��H��k�{���_DL��~uL�B�7������m,"YL��t�=ῳF�F����a�X�X�r����}�D�w�����%l�w���y��9.x�vWVrpeh�F�`���{6��\�ED��,tX�g�?��oGͿD�\��AR
��$�����ø{���k8�J_�rJj�iU�mc��;T)����[��}�욈	/�����@,&o��� =�_�!E",��b�o�q�����0�3ΪyK	�l�ţ1��vǆ�;q|#	��0܇�������.����έ��3r��9v��=�
��^�T�~Yo�����������q��`�V�b�BZ��)�z��w��x��'J'��^JS;�;�7C�$�,#M�:@t��^�a1o]T�چm�����x����n�=ȝL��t�F�y����f�ޣ9���vlAM�¡�#D�`#�;ډ9}s�pw���P�A ��3���82����i�o2uG�>s�A��
L�U������LC��;TP��9q��S	�.m$FV��K3ĬnƷH�_C+X�QW�'��V��M�hGw�Y��*�W����o��rs�	�\�O�C�	[Ux����ڼN���v��������?�t��ZT̈́����k��ZZD�>��"j"_@d?H����m�*�H6��mF��g��9��0�p��T�[�Нڎ�g��S �� �i�wڹyQx,(k�9���1�[]k w�
K%&�u�ɰ�U8�'�&UPȟ��G��fr��("?V�0�T��K��Up3���}�z�e�K�٥�_~��D���|�б�/4X��k�F�	��i�ϒ����1k�,uQ��pq�Te)-���N��n����Lh�R���3���.�0_KͿ �,��çS.pr�n`Y��J�%>�.dm>��2/��l��V4i�j��Bޠ�w���xg�c����"0O~a��"K�<�Ex�VZ�����L52*]��|V�%�OY���A��
�r�Yѵ���%���p}[O`m��< �ya����/Z9%�103���w��{�?�슫(�h�P�!Ͷ�d	b�W	�8�5��`7mPY�����2���R�\��<t�O�d�~,7BC��WY8�g'�3����Z)��;�29�1�2�ϟ�[fLm�������ܘ������4|:v+?��'~��zw��.�ۼWHt�d�.Ϲ�� ���������'e ���{����eZ��	�A������d�S#?C �ԣ��)� 4�8�5Nۄ)i=Us8���u�>���	�y�:���b�*�]E���qY����.ZUbd����J�e@@��E�ݘ9Q
��-�@�;1��Lu�x5o���nP{�V{�<y_�LeU�"�,'��s��2[�4�� ��Jb����mn*����s|;&P}���bh���
��G,I��G�����W�v��#+�U0	x�g�����
��X�N������"Ɖd�ۑ�"��i �Z� 4��J�P:����e곛�v�SX/�CN��w/z E���\s`�C��Mq���v�c~zv��;l*�P�A�)��+m���z��C�Wts�N�Z�	��M���	�r��x���G�(K���z|]�"%� T�B��ڢj	���ٻ�����u��%ƣ����@�T0 >}�F��PͶr�e���0yq�ӝ��ta��h�{8ݔ��	�:Z�_[lt�R��b������&�K�)/��3�}v���L��W^[M���%�]�|=�?���K������o�\��3��/���`ӱ�ϰ[���������"�X�2��9G��l�?P�]�	hD>����b���`��a�M�t�	�TR#*��x<��#cI�Llj�$����z��1�&V�}"�oxE�c�aJa�ż0����>3��nK��߳.S�hRx��F��@Y~n�9���B���v@g	���/C-��Q%��b����-�u��o ��y��x���zيX|��e�0nMk�a1�r�t#�k��������a�ȣi�Y�V&P�Y�
��vJ+v��&R�K�w�r��� �km������:^�t�� ��^���E7/'�F_S���:�Y/B7��՝/�I}��g]�ה����x�jwX��q��aЩq<J�Dm�Ex���uNwP�*J���z�LpM	:��_'����ߝ¦��w�p��ݦ�պ�ݢ��ĳ�����E:r7��_��Kl����@r����}�،9��8����u
���f/a2���'a�E7ڻM�m��6lXJ/�>t���a؉П���4��t>��_�2�@G��=�H��bs�)�����Ea���dJ�҈YN��j����%-�TB̪�3Ʀ���n��M� ��[l9��K��§S�(3�x���xȜ�"�KT4�!|؅�߉�L���G���#�I����9�=��=P�)���0��p�5�Z%���m+� pu���}�����I��`���%*�[0_�Gq�|cZ?]�s� ��B`Cn�`����a=�T�B/5A:�l�З�)ϖ���
-��J\�e]��/Y͵ߋ����R�)����^|v8n��6g�睲�7���iv���<�q�q���'�w�^�t�=~��0����G&S�i�ê�7#����N	��LkW��w�#+ּ�b�ZD�@X$^?�f�f�O`R=��F��L5��P�& ,MgU����Ȕ��`ӫ+�Q��4Jj�*��J�L\�3�Jl�5mx�Gd�ˀ��6٫t�qv��0�'�-jE��A�J$c.��߄gFy׼��Jw����ܷ��/��W��&i�	R���H^AA��Y��s���f�?��� 9+\��P��Y�}㐠2�dt��u���s�'���=�Ft�u�u�-G9�֧�-��:�d˥�<��8��h�2�tE��<��"��795��2�9�#ƍ�伢���;��Dgν��ɨ>澸2ʀ��2����	^���p���h�W�`" E�t�ooq�=w��(,ˍ4W���"���u�W�8$�����Z�T�� urb��Հ2}��SEF"	��`�0�zlO�z'Żݣѣ�-�$8��j`e�,�9k
2ɞ>�
1�(}yW0M����Bb���ͯR��J\��}�[�@V���u���H*�x$�d3��`�EH*Fz�.���e���J��@ѻ��ߜ�H;7�/���[�N�'���@�v�ؐ��p�s���2zbE՟b��F��k��{�	��a|�X8�	��5��ut�nseYP�Z.�I7TXV�xrI)������9�u;T@9y��l�RHnQ�1a���%�$�Z�ފwZ��@O��D�{��x���Ja��SjI�y��>e`�0���G��PO�&��$���L%]�[N*|"�Њ'�E�(�)��z��[.ʒ�=��b�����HV6-,)�N���xSW��Y��[�5�M���_�ǭ������n�~���bd���X�����t��3-۵T=$��U�j�Q�>��J�F(��I�a}g��U.�	�H�������u�����!��F��]�$����g��Ki��[����՟�����r��'T�i� �z�b�ES����1@La]O<tVG���^��X��2'�ў���ҿ��seX�A�x�8�Y�u��~�%�Ⱦ�,�u�('5	�J���ڛ��I�n�sdEW��5+���:��ӹr �f�8�]-�����xyC�:l��� Y+I��7u|ɬvJ�|�� �V���fv�t/����������.�E�C��:� �b��,��CP]C(F;��
43F{�߭�;��p�ݞ'Ic��`<�Qsh�dO
`F�I����Si����Q�=�ay�ȷ˶:����4y,�Β�z�f1�z��8�*�X�ʙ�"�v�Sf��5׭x9g痟[��!��r@�K���N}���J�<���/����xg�|y"�:!#
G%��`w����d$�%�4,���:��b��{tU��.&dH;gQ,Ӷʳ�����dZ=����i�U���tI�����ϻSv2v�<�����m%����(h9�"��Ej�@�=�| �q��e�~�e�@�0�_UK��7)��;��-�[IK��;���}+��{+�v�_�5��P��)�V��cܗ��q���I|4E�{��'��9G���2>U�e�g�����4N�S�+4����������4981�S?ϼbI��
d	~"�K(��g��`=��[E��S5�-��3��wS��hi�5��2U��&J�IE9��x.�x�����]6z]L���qq��'�A��N��hҘ�Y4v��K�E�!X
�i暱�����t!���ڍUZ�Xb~�š�̷�_�~@�cGN:lq$!i�j����@0F�OK��2F�c�,���?4��Rp���tM�׮�?���m��>u����1 ͳadaO���R?A������9Y4r2�/7_3f�nj�7d�{���"�h/р`|
QeN0@�l���4�����|�8�Vu������j�ĉ��-9���Z�Z��N��?D�������t>�
 d̑�,d`e��.cqȤ��X}�<	�E���5�8QYs}	�.��suSqUn�S7x�r����%# ��I���톟pN��yZ������Z4�f��υ^yz�_X��@��X���L-�Uo�a�h�1�����N���T!��C�
o��ɈcL Z��3�f��=�
�l�h��F%�ߟ�˻�3oL{�6<��1�ap�qK�ʒ�����$���v��B�Ge�1��C��W��?�aEW�����(>iR��q@�s�B7�ݗ<)+��| S���l,�$C��I��NG\������S��� è�5m�t�V[u;�eZ�ُZtn�H^N;k��C��`�^ko��J�]V���ȁw�Y5N��73��JC�������Lq�ԟdMh�$ƇF��rQ�z���S�M>4i��ߌ�@%� 
V�;d0������u@|uo|^d�
jV變ߎ�Z���u֩�];K��>��)���?�4��ֲ�O�i�����eÃ8me#W]~��N��!Ԍ����L0B5:m F>�'g ��Qq��F!�=�ܗe=� jrT���tʅp�l�9�&R��������  �b����Hx�3�����H�c�K˫���2�2s�����q��́�G>B��M���B֎���`�(I�Q�	��݁0@ N�*�6�76�[��F��R.rA����L�Ez�1������wl�;6~��Յ(_Xp��w��^ѣ�B�
%{�KF�h�D�z�3öҤr�B�^Fi�/A��ɤ�I�܉Ӧ����yΠ{*�ό��#��kP���S�i�D F�
Ye13���fJ�]��cJ:]�x�i�~��R4�26��]�;�ĢY���nL�^ky�o�e�w\t|���z�B�T�V�6T�J`|�v����^�2��ȟ[��NM�2�j0f\�G_����۝*�;�����|�ý�"�R�2�"����8Α�4;��H��;W'�pS�%XPb*�@3��!e�s��(h�PP�"P��}]�R���"=15Ģx�-J�]�����$�G䈰�I��82�T"���~��cN�lAE�2C����(��!_�T�>D���{e����|r'L�i���8Y�?!��&'+g��uH�r��p�`��$�n�����z�J�tB�{b�yb�vd�f��B^p��1��⢶��z�Cgi+ny��5ͼ����j:8�O7��R�<�r"WG�Z��2�{hѹ�
�0�y�b��8����rXRZ�Q$Z}F���&�f`o�F&�}z�k�0w�>�s�J�	.���u��K��s c�$�jh�u6N9�8X�8�������m��!dw},B5�׫`������#N�q����d�Dh3}�� x�F�%_ �2Ƣg��-j���ťGϕ��=��#b4�c{��x1Ϭ��9�Et_�`�����苍�q8�f?
�RF�ap�r�5H.���f����H.ݒ�H�!N���΅����l!Ҍ���e?��Q lt���iC	����Ad�B�𒹞&�=dl��ۗ�T�2�'Hg+�����<��*lF�Djqo*W,=zZ��.�l�6�f��Z;dUd��8� ���-�ʣ�o8�1�L�v�8-vN����&-+�Ͻ�*�9�\ɮ��
>��p��ɕ��I�ZV#�b����|!Q"��D�ܙ���=�i�N9k,�ի-'ܟp]_'�U����MW�wT�����΃�ȮFQ�PX5���~鳞A+Q��g݇ Lٜ��4���!.z(����e_�.�F�0fڠ}5�U+�+G�R�/� �_���Sm��XK t4%Y���k#3���V��i��"�BF\Y@��˘���=I��tQ�%m�aOG�Lx��r"z-!����xRmc�V��#-kYz�l{lC���� �5���-�:Мf���a�#W�ᗩ=��f	� %$nm�YW�k�w��9�!ڝ����{6�H~7�^������.3ֶ�������5�w���)F��vࡐ���]\���Ɨũ��-F�P ���a�mZ��ٮ
�����&(��04�	��n�L�b�����as�eZ��o]�S,�8i��#��k���ꎩ�Z��m�cS��{�Sb�w�>��P������7ӭ U�i�j	��H-�~֕���l�p�������L0�)S`�=��\7j,_�6P^=w��綷�7A��s�fz� x�k� �6����x����y���%�u����%o���f#�d+T�j�����>�!Ɛ��4o�3�6�� %��Z\p��rC�$@� ^$�;��GՉ�T��VI5�р����罼�^S�6�g7j��[�h ՜|ljONn@T:��#��S˽y'"hk�2��iG��gڭ��:m�,s�%lv��#��ܑ���4-�o7�2�{ ��U���Tm���;�c��Rɲ�f!i�!�i��(��ֹ8k�ᓲt�.tb�_�d0�E���MƜ�2D���������t�L�p#��ú�Fo���'����ބHש���M�B��6�]��E�+��Ɛ�Q�m߁�MC���2]��dr������R�L�7pi�Wi���'���CfPSw}��cU��UD+��4� ���f ٬g�l6�Ly���y�T�v8�?�`��r�˄��H���������N�\�_C"fb������G��w2�봑�
t�8K��4�oO�#W��g_¶�ƺ����|6���4�W��pV�zC�)�8�'�L�fbF�y�g� ���-@�\�pH��F�'b���b.�k��N�����/�%�-Q\Uz���Z'P�uRÓ��2�$8�S[��0B��\����������VY��}�g�Ԁz*���/ƭ�lz�'�����j5IV�FR�^$���ߞӞi	ɻ)���N㉴�P�{��9�R���B��Jq�Q[�k,#F�����v�4A8��0�߬7��!��u0��"���t��h�ܪb
��X�8�D���W�j�Bˬ�wG��S\O��]W!4m0^����!�ԋ%�U���"�r��R����sY��~��Y,���Q����6���-�O����l�"�"k�=j�y�;�2�{�vf\?ASi��S]UY���u���۴���0(0��]�5���i�����@����wnP��������鿐���Ә�ڼ�Ƚ5c�a����B��\���eE ��6�!��/��`3�S�
�G2A.I��:?�V%�hk�W.�NtT;��tQ�o�4	� t/	o=���2eM���h����\���Y�e<,��[��$���&Z	�|<h�7b����|LSYAhS�@o�˵Ñ�VBm�yɐ��0�������G9����r�	�*)�q�8Ó+j�W��#�=��"PŎsϼ���i���v<�!����O��G�Y��N4���"�Ԕ�F[�;�.��J + ���� ����0b<�D��XlxV64EB    fa00    2650RC��`�n���?�`펫9FG���$�#�2�a���h�aOޝ�9��sM���� J\Bj6����M�K�o�Ai�3��'V��Svz�� y
�H�qW���֩Q�4vv{�l~ų|8�j@�2���yE	��[hR#�tҳ����'�}+��fR:��}|8Oq�5פ��r�jP��dq�l٤��臕���(׌f�0���Or�GS��TTIQ&���mI�s����Ï�������5�ѩc2����DRL,dKy��NE]��^�MlE��Mwl�N�ڞj�J��� 7���ee�EJ�/�����Ά/d��^a��[�S ��F�C�04�nZ��YO�_��}{3�vĜ�\)tƏk|�����01%�6"f�qK�]N�)�;�#��NZ6R+dݒ�=R}ҧ?՟�C���
������T�O���@X;�H�h�jL����7x�1t��=������o�R����Ҁ��Pθ,H&�w8�!xWR�(���l�'�Y��.�)�E<<)���4Krr��YôP{Z	����)"'��e��:;�-���\�<���k��� u�J�҂.�Yuk��6l=ü�p��Z O3�o@�t�Vj�`�b?�� $1�~��r+��R����	~0� ����|�G׬,X�pοL��(G�7��oT��C3�^wP�y
�e��âM����6�&D{:s[�H%o[4�YyU�������R���`P�I�;�#z)�K�����^��#�+��$�|s�������nO �
�qϜ�V!�u��z�˄�,gK���۾,w��S�)1�B���J��m1 �=�d$��l�m:ӧ�+����g\�(ZcW�
���o��ס �g_�L29s���U�O�OZ(Ew��"���a-uȊB�ΙV[\��5BS���ݖ6�)m*�6�2�Ea���4��fc����:JN�!��9PQmM%��G��\F���ӓ�D�m�.Hp���b����my5�Fw-5�_�ˠ���!`�V���0&Rw%n6֖��^ύ���L�����-[F�����a�c�����8A8#[5�f���X����r(*�S[9�<nG�Nx�zTU���,]�V�"5${�:��Y��X}���.̉&�iȄV\���AĄ��t��2�<��hk�\ɾ�{�*Tε�W�{���<���z1��Z��_����ӛ<� 6�-��������/��� ����Ċ�� ���N-h�q°��ۺr�V����h*^�e�4X�r�+�P��\�}��<��]u
����db�.���;��(�5�)B��іg�0ӉmR��M�:����[�C����Mi!*/!�仔��6���l�~}q�'<��R��nF�/�9$8z�3���U	w&�\�ٷ�Z��~���m��b�²�x�w�hD����$_ � ��5F�h��!q5��չ����6�Qԫ@ip,;`GT����NB%O��+�Lqp���x�3��[v������S@[�=�LE:Q��F��o�D�<Q���'M�����վ�~d X��OWz��R0/6f`j����w���Ht������af�y����H��܋�h��������M���~'Ȼ�.8WD��[h�R��A���eFH#NEz��m�Ve�Eؿ�No}�{g�{"�#S����O���a �vUQ.}S��8A�Ӯ.���b��[K-s	�����z�4! !10{#��L�1[T*��}_E��q�@��+p����1L]�k�Qv���b���vI5pf�z�� �T����	�vѣx��8T,�y��<��{W�e�|H�Z��R���%��Gɜ�f]<k���Fe����������f�����#}��Yǚw�`ru��Wbc?᫆r ?��g�g����L����'h�@��?�3���5T�u�X�?�
�{�����f��,q�����}4R�7_�^y�Z�ة�~�V
r�>g�\s`�����)�9���i���=��ho������Y��p�s�W�A\�@���#"r6�r��R�H6pmO&%���K{XsXkU"^F��Y�����(Y,���5ԿX�΄C�{�g.��Z����dp����r{\x﫽jD��fhM>z��R�7�����KQF@`r .��Lv*��ƛD˓Ǭ;V4 C�6E{pь�瑃����J�e�����A�Al�lJ4�J]�����]f��%H@N���������v}����q����cS��������$^-V�-�!�����i��@����zu�И�5g������d:�S�\F���n$Z7��G`�R[��)P0�r�Y�(���2��1�k�"�%�%��c�������v�k������ �j �et#7�j�,��Q-�z�c�J��� $����^Nf2�%�u��-�����O$�6i�*�߀9 �՜�2	̔�ϻ�����s�Ed�L\X��}%eCQ���IXL����@�6�������P��$�&9V�Cғ��C�}�KSA<* ��C(U����}s�(w�IP/*q�x�;E_�P�����69�k�XF;gS��>l`�E��ԍ�s{��M�n�y�vY6~M�N��m��}K��}
�I��e��%f��S��YǊ��\D��Ĩ�	V�(����}��	4ņ�W�]󨸩
�8�E��aqs���Hw@!�&�uh�	���8=��o��5�̪�A���U�a���6!s��@��Q�"l�d�6�ٹ��7�$�X�UK�s�'K�w >����Rf�x�n�6������v��UG
j��FP�G�U��?�U������{��Ň�/E�%p9�.G�{?Y�|�Y�0�h��[�cZ/cW�
�ey5CA*����j�dd@�/�vK���2H/�(��2�g,���8U>#3�L_�y�ֈ��}�K�Xk<�NK�/:����ZM)����K�Q�	��h�$\H}'T���(@���9J���a$�$������ �6�.��k����wW%4�9L.�ƃ���8�1��&���ɐA��Ǒ%_PB���G�6'�U-��ĬH����0�FP>�(2_mNs��[�t�&f{ϗ��΅���'�f.h�D˔?�,m"����N��pf�=�"�\�1��~�w�/�v@I+�k3�K/�Ύ1��]��wnj�dF��'
�D7�j�y=�~���QH�w�P�`����>���0m�/��_H:�{[�r�r��v��q�#��4�KJ+���\��s�������5ʥ�a�ʢ�����H4q�?7�Ჹ�`�����ay��뀿$^�a��h��yӠ�D|����O��P�O@1��礳���k�]�Br���-2qʆ �H�iR3!���7�{ˊ�?EK���3*�#�.��"���8,�>@���.�����X?D�r�=iD�ћ,�KYJ ���5b���dm��h��K��M~aB�3��W����h��w1�������Q�Z��w��=�4�Adto7�$iI0�&^�f�%�Dh�E8N�E���H�҈�0�P0��?��n�&�E�k��2�g��g^�t.\;ݦ! l�X�c9
���9�W��By��l�;8\�r}��Z��ޗ#�M♨���4%vn@����v8�n�hƯv��j m�	
CvH?�sNa�Ns1cɬ�{�������(7Ӫ��\s���B�e�4�v��#?P̠�����º�������'�錷�oFv���%�hS�=�ܴ�r@r��6�+�{�h���h㼎���K��g��z�ۨ��F�E�5%��tcX���ʥ~;��0��b%h[K1]'���@�FE�c{4�o!"Ms�l�*��Y��5jw,Q�.S����_[q[&{�*���X�}�a���.���2�P�XKm��ʹ
˔Ϟ�A��xߦ[p��o]�?GBw�(���r�6|�m��۩ҕ�u�S��8DU3^��9�?h� ��g�hr�m�$���T)�dyw�;m���z����;F�Tyf�}v�s?ֹ��K�1T̖<=����B�uL��q39���c&�>[�����v�W!܄���I��==�#g��m绀Ӌ J`��ܵ��'6ڳm9Z?h�^q`B�A!���2���WBx�z��ck�f[��L |=��B�!x���[p�6lt�ޏT���������M'ո��ʹ��Z�@�R��o�G��}գe i��[�첷)����F��q.�-�s��C���íR��}�
Y��L;O�� ��TBD&ƫ
���b3N>J�K�����}�t�AFq�\z������U�������{��1�r��O�'eߩͭ��WɢR�k5�F-	f���F�5E�I���X��2U�Tv��ا7mе_��d��B!� .���'�8��J�{�*G�M����-������	��S���˥p�L�t
�gկ����x��]B��9u��z.D�U:��*�9B4^ ����w�a���|!�5����"�����Cd}m�(�6���I�9n�nۣ���pt�M�i�{6�!�Ou��b3�J�~�Q~��W0���/����xq���#�2���r��e{�PhN��	��,�P)�Su��@l���w�O��%�T�^�{ ��u����,��EZ�k���t[�v��z��֕c��;d�y���}G+2^�X�;L��ǅ�MN/Im/���w��BT�O�k���&׳����Vwi���s<��y���zq���|��X���mʅ���RP1nby3������d�	�V�!C�q�:�Q��Wt$o֐;	V�Q�+���Ӷj-|u�Pd���A��&���k����i ����Q*�������sC3X��Lm�Ko!����>f�7.2����#�8m{p�������7��?��(ߟ� �P	dM�\�������Q|�x�/Ua<	���aqp)*�%�ʿ��@C��G���O��߂Q�2��K�WR��=}��]��%���6TS"7wOq�9�V+x�TA�g�,��}���|�}$�.λ��At�~�zD3U b~ö��cp%-mD
�tS0z;/���������T�Λp"�	�X�81�8���I��l��o"s���
�u�ة�d�iD~'����:�B1G��EZ���6�lÒ�������)L\�[��ڑ�z�W�$�+�\c���r�"t��P{-��LwԔ�kʈ�>�L�lb+�DٹZ@���B��Ή܎%k�����(6h��0���w��J��_נ[qg���d�wRR�g,TcO{\e�����7��ōm����8!��/t�v�Hi+�>�ސ��M'x��JĞ�o
'�)c-��#�E�h���1�se4�����5l\0CU�GM]'ɹ� W�/�A����R2Fp��m�Vɰ_�0{�\���hU=ȏ(��@�մO�5q�}[�v����<��>T��0�w%�]�rA�w���}{l1(媤��W�~�����F���6�:ۄ4��-�W�>eR, x���>|C�����2�+�<��������wk�M_嬒'hvo��\#]r;9�NGPV��ul{݀8{�X����7��������Tu�5�@�Z�#jG�̄�R)A�{ Uˮ��f�?,����`�'��E���9�G*N|U��x���;�m�N���.M�4�3�������L�:�ռ�_�>��^�'���$�7$����*`ɢO�O�,����):=�HQ��V>{̕����@��C��&��"��M�_Ƕ*7	��&����U�� <�hb��b�b��o2���%��\ ^r%$��[߀�ic�N,Y���A�bh�Q�]L���k��#e�9 cU�RT�����a�o6�=%!9�_pe��pxc�w#JIu���ޞ���{�)�U
̝x�f�t\(rT���/$�i�P!�JI�����ÿ�lw�]����g�Ci}�����'��W�k>S_1�g�I�2�	����`��ҕ�����^���	��Ῠ@f����ʷ,��Qo./f�(��M���y.;u�t��Q�7�U��I��D�E+�X]fF1ŎR�qP>f�}u���_�f���TӤzp��r֘�:�Su��@���c�c��>�W
F4��ή��&mȰ,Ӈ(��)���)�|W�M:z��D�K���ե��R�>=��[�oڲnd>����.��]�������}O�k�r�'9�]��Pp���b�h���蓩8���Le%g&��Dxo��"J��O�Q|x+�LՔ�������x����x�| AͩƉ�� >��R���1�6K�;�����¿M�m����
tۃ�/�h)��ŻKlD�O#=k��@ ݛy~Ӯ��.�YgXڒ��Bl��� <mc�l��e���j�݅��G���h�'�R�x}����9I����_�}��4����	��ǧU�;{�`���K]�+fw�0"���\���"��/��̠�f�Z���ղ$0�(3H �+W[W��F��X��Yd�^K�G���Ķȿ%���s�O5���,�������b+�8��u�����7'�B�|j���2�Vެ0�k���S������ir���Zך��,��@=>�.( ��C$�4e�'�nj�`�r��5 �4�ڭ1F$�d�ޥ5�T����}Wn?�ڊ������<�p,�_S��)��W4���8�z��-��g���V;��\NoJ /k��Nd�Oo>"�J��PRme-꺁� �fI�S�r1�
z��dU#rl�Z�"�5U������<���+�E�*��NS��[�d_y Rly���Ñ�ƒ��0�<�2C7�	�w�� �a�l��ZA���ib\�A�Y/����["�H:{i-��8���B��}��$<������-?�~b�o��D�$U��_��܀�*�Q�l�*~�?�Ϻ�h2TJ������vȘΓ}ǁ�TE�=��H��P��Ê�����`>�R����k��?��l�uk�#uE88cR��T�wl�	����\�ꪋm	�*��55WT������l��H��ΐ��f��+�\~ k=�]�bW�dOZ��J�-���
MA8�����ַ���%p_G���̓bj����YP��O�DhܤD�X]`���ḣ��("ĨH�9o^�]W�P(��a���p��|.��7g.+���s�<��'>�T=ݸ+�л�`Gs��,W�i�n_�c��;M�`��(~|W6:l�x��@(�K�dA}p�n6r����	�*L�Xku�Nݩ������ݺZP:��?��='��T��ws��!�8r)s�kX+t��pd{��>4!_�^��9�5
����h�oO�X�Ҭ�؞9��y�9%Q�.�x;'f҈%�v�;�z檡%�����3&3�P'��p=%�ִ���j�ޒb���QԘ�S"OI���˅��le��e��:���2�8B�����d�N���v���V�"Gq���`�^#��������%��M�I��Y���D^ӗ��o�~&]*��#+�t��l�ˤC�aTJ���<^����B44�'��'�e"��	=�R�r��qa��v,��AѰ�9 ��N�_׊=��L�s�~�����5<b2��W�����������65�X4��7�H�\7�[H�Mǰ8����f*��_1���ex�?���s9�A�P���a�*Y�£Hryl�����a��N����]Ö�s�`���A-�V��9��JN�N+ȥ^��Q\8x���������jzOEcf����s��>7r��}k�tbB�S���%�R�C�"�2mI�g� �A�R����v����MoK�<���Dv�����V�k�,K}/̲��f>�����T�{�h�(I��C��A��Լ,EBп��\�Z7g��%���U���8k-Z4�"j5�2��o����wij1	mխ���P���Q�U�A7mU h�&�j��K���綪c��x����J�=��~��tQ}���p�ӓg�J/]bʏ2�O�Ba�g�<&b�cy�׿���bp�r�Ӫ��c/���#qI�Cy���q6�b�4�4��u�W�<��Q�s{���S�)e��h���<u����0G(��8ko��FvV0�U�0#��V�,ă`�cʼ���Ñ��+������韖���d>�42cCo����,)�d���c`"�Z?������]���I�%�$�����?���y7g���X0�����G(����$%N&���|�#�Ƈ>t��%7cGA�k�b��������^�Ls��I��z�C����+B&�����I��� �j4cCU���z����ڇ�|�b�X�J
��8�B���D�2��'����s�(UE�44^��@Z}&m�t塖L�oDU]+x����6�HA�y+��\�$|}���|I���w�����΄�̄z���I�(dlہ�����0AY�a}İ+t��-��k�D����߾�6Xǁ>�=V�'9��گ}&�L��.�,���moe��Q�U��sZ�1`ibs���_C�G��R����u�?^4Hփp��q�t����fc�?�d�g �DX���h��Q���4r$�aF�'#O|�����r��P0@���|�3
���wh6��ƻǾ���҅nl:_DT�-T���1:g*+�)����O;xB�s!BB�� ��Ǩ��aϚ��:�3�����CY��=�l=�I��t��Û�X2q���{�ɭ�Y!�=+"z-l����e��`��a*�2��R�T�\�/���`3A��;����$��P�j8��&�\Ý������+ؠ�.,��E���'�����>f��5ƍ��񄐉�}࿂\�춄��B5;�?i�4C��L⚞	����2눳���o:9��({/Ͷ#1a��!��yd�3���;nU_RQ�EaC��ҩгv��F�T���S��/��ס��/H�����{����|l�r�U���}aB�~.s�4i�jB�LB0�k�q�c�p�B��l	K=_��6�=�E.��r��[O�h��c��\d��L�*=Ll�zN��/YE�j8z�\�_��ڸ d�
�k:�q%K���P2C� I�ںp�o���N�w�ւ�v�gi&����������:ߣ5D�:eJ����2*!G�c���8��w�R����I��WH�c0��E�	����b�sXL}I7
�8'h�	/���j���6N���p�����A����7���)䠊���C�~�_�n�M�ف��Y/M
�V)]��0��ۗW�9>`�? qӱJ;-�%\@e�J|(�� k�y��sv�^"��l�)��f�QM/ 3�=2�y��ES�6n�����r�:��_�lU���c����# ��h��`~+����X� �(��?OjS]]H5���^%�Di����dN�^ &-f̹��e�����w�rz������� t�*�]H[!]�t�lu�d�	��C2\lur�>�ؽ0E��|Yu@SF�I��F��Hap�i��|!�&6������烹 [ɚ�U��5��c���m��x;���:�ە��H0XlxV64EB    fa00    26a0����蓛�x\%=;� X��D�S��}A�a��Q:�W4�8�}�E�?����ϻ5x^��훎c�0���_ɏP[[1�����㐣��X��|�#��d�3�gχ�&�jn�o�Ý*=·�4,#f�	/�J�PIQq�/��<M�$M��]��B]�)X����d}h�.����^"���2�����)��f����ω��Vֺ\F�'�C�4���d�Ϸ�lr�ܵ,����^(�i�r�՘������[��*d�=N�EßW�vl�y��6�0�_�`���:���!E�)��w����ߩ+��̼B���G$K�S_G���{�f-�s+p,3�Y�c����O�1�� �;=D�h+�큇�6z���zi�њ
����V�-׭��K��-���Y���"����/O�/ͻ���ݗ��(ީ�^]ǣ��?���3�,zv١�ၻ�0�v����{�)"���9�'���n���S9:O&��"��2ro�P�m>�ȇ7~ًO�m���p��WǇF���ب��f���%1@Z�e
.1�XLW?���>K�I�E�Fmg�3�w֦�"�\��eѻٱ�#�1���>c_9�Yr�QU�Ù�po��a����i??)V�Y� ��s����7���`�e<�x����K�Y��[=�Eל�Z0�}exfe&�`��Ƕ"b�����_�F�5䧍�=����4Bc���Y7�|Z��EѾptW�����%�_a��0�Y(=ae_�xLӏ'�?i������ޖ<�߂D.�|�Q�~�����L����B���mlYs�[u�̵ �KO��%ib��P*�վ��ٞ��-~ �ܑ�.��x5�����QV��e���[�r�=KM]�����[ h%U�f�ϒ�?�?��!*�W��~*M4�[f�I7G`�hV�3NQ���4m1�nԪ�P�����_\����vH��<��9��ڮl��}'�u:�|a��IF3I�~����&���}�ݪA�;��Q�wȝ��+hmVf�S�;��{��^�43P�����~�s�;ᶼm�o��7k�"��k�*���Q�OxmG{]SLl��w�S�w�F�3����}E�Nؓ��r�۰��� ���n:�����%�?��<0�u�+#K���2n��#Ji5�۞�Sr��?��
����g{�ǕVJX��Tȸ\��0���`�ro�;6D��T�mIvj��qU��y$et�/`(���������b�����ә������@t>�"%�2X`;��Gr�z_;��mMђ���8߮�;�>p����u?��A�h���+��+�-��p�h��uݐ��xA2FaPr;��}���5ڼ�� u���<�]�,�N����ZH�߀-6;҆��K����z+��V���;"L1X� ���
�g:|5'Ա�]�ѷ�橶�vg&ҩ��vL�b���a{�ʧ�%�����p�喇����[�.{�y���i�>
L,�6�&� �	��qZ򜉉-�-�]p��d4�GA�Yc�#��nz�-D�﷟x���%����_Z%���^a����mL�:[�g�990� �x~�"���L�
P� �=����!����y|4I���9W}Ԇ��)�΋��w`9d~]�u�B��I�v&)� /7:��H�Wc�����N��U�X6aϳ��?�'7O�MT��ds���{Q�P�$�N�Z���gLgby������_@HШZ-��b&�(VT��
��&�]�����/�K5���Bd�����
z�L=U`].�j`]̥�&�`�xm�������"��ebvPoh��d���]����w/�U�&��].�1S��pҁa���6ڊ�C�4mse T��Yu�k��Sξ�KH �8��4�?�2���uc���*(/P�[��V�=�xɼtd�~�X�|����ԣ4yr8ѻ�-?��L��! gdMJ�V�B���G�J8�TΕ�Wh�P[ό����/�a��n��r�vX�g��d61O�����t<N�k=j�ͨ���?��>�[N�5��'-R�n�Mi+�=^'L�S+uF�$�mm-� ��ZTɶ�,�޹���F�!z�8���x_IL	n S��FA 2�}U衪yT���/(>w����|�� NI��+������<����첍�޶Q�$%�ݤ·rm�!��h ��R�h�ɳ0��ln?K۹���!*TV��.9�}~�6=0ԧ'#3IU����ǜ���v"jO���Fn��o��r�.��B��T����ݩ~h9ۣ�������T��V71��ZeH�Z4_5-�tf��V����C��cU��YO���D9 j.C��@^�t�^m8v�N4H3���c�<�g�����-��<*��{qЫ�Η��8^YDƖ�F�����X��^��8s9�g�U2�g�埢�
}ms���gv��*�Q���=�`䫺�+�R�LT'w�å��Ti�p��;�����ϥ�$�=����IX��fQ�T
�r 2�l��ՠ�/���E�?�fd���K���|/ ���(9���j����p�Z� ��J&�2�G�݊�Qm\b� �!q�!�/`�ȭi�֨B۳-����3C�>A��-͹��u��) ��[��:��(,�s��#6��ŗ����$�����?�93�#B^�GF�����q�/�nElO�ݍ�6�����x̐�N�%�V����Q�H���ȅ��X��Ɗ!;M:�OK�j2K��}�&�.e(H�JA��u�(�܍���M!��Nv��^k߿���'p����>Ĉ�Z8�҂Go���9D*),j��c\w�� ��t�	S�3��kSCU�:�&TUE߳�:��RY@��`.�X��h�S����;`=����߆; �7��z���ƨ���2ew��J�+B̫=�\B��:�_��ϒ�lj�}�����%H�* 3�`���4�'��4������ժ}'�a[��M���ǵ��4C�:U㧌��ӕa�����u��\�dQ��t kꛋk���e�NO��A4`��nA�D��qϭ���5�B��W׷�k�FN�f6k� �T+�|}?�A��.|6?dJ7 ߝ�ci�2.ŕ�q��b�ϴNB�t�m��o�z�8W�i;�> �M�q�~Z�*r��Twsp�oo$��)����*Ae|2����6�S�J�e�y?�s��1�/ǌ���O�M�:X��wC&���9��^��}��˩�D\�
b��8L�A2%-<_'���g��d�`�����H�I�D�����|�qH�y�Y!���)R�' �d[��+	��=猙٤����ra�܃�p}�Q��w��V �?�Ys�n��y��/0i��@�y]R����N���R�D++�&.%ѫ$��W;Uu��z�n1~Z�rV���	7zXYLN侉ׄe�����g�g�#ح,����;{�Z0M�>1S[�?��~���W�;��S�^b��"j�8nwD�ʨu�[ �*�z�^O�ќ��WC~)qB� 4���.k��8Y9e�E?c�|�c�a����F���֧�G{�ਓ�,� p_Ϸ����q�9��x���Mг!A���P�|��@�ox!q�d�j<�u��|ZC�[�E/��,hS���/��G�V6�E�,z0��f�`�J��I��"@��Ü��d8�e��a�fA\��ylnn''_#��j�E��)ċ��- �]ou�.�7D�k�K��P����BH��{��d &^�	��׆U��15�.�%`�3�D���b�8N���G�0]`�ɜ�%C�	�F����p���	%�&�Q�̸��H��O�T��xͨ�]�4�PĒ��ׂ �Q���F~�m=����3��<����>�e9���g2 I��� T�QF%���<�D%T���Y·}e%�b�hc�.�ԵB�K_��	�⇽wU���ױ ��\`�D~�a;;�#R|���=�Z{F/��'�� ���&1�	Z�wl��܍|����9���d�)i����ԏY[9@T�o��Zg�(}"�����[�ۺ	��3E�WN�$���rD��Ɖ����?k���[�������+A]T֯)�^hf�.
� {Xւ��U%Xf�ho�F���Ҥ��bw�MR�;���w�Q\�::�2d�ƻ��r�:\U�o��ڱg�t_� @���L�-1sEX�^;�O��=��4�T�mJW)e�2Vv_]�~�A@R��ZsѦ�VV2G)F*YQ�b��$:Q���F�_!ӂ�~}*(�[uB��Ѹs�A�����;��Ŗq?�6��oKI��k-j��<��Bx΀��p�/�I��j@�)��� η�Va�"�[cyS/��`W2"	����4\b�30k��4_B�H1��xP���D������ʿW�5��k�	��������P4Dh�=�\l��a+2c�î�O���#��(��#ǖ+]8U7�������(�\C��G�)��Q��Q�w���p�,�< �O�y�ޚ���
��RR9�;�n+�g�F[# ��쌃��	g��9fc
��࿽�b�	(��ِ�C3M��#����N>O�V,���{h4�����쐺(�`�j��P�G�{�g��J�A�Q�3��
��M��o|Ҷ�M� �k�_b[�uP��_B��@l7S�@���-s9G#ɰ|c���&xT*^�(���xd�Ce��vM��<�H-V��/;,u{�AKŶCI
�Y���c�^i�7�sUV�7[U�t{��(i�h���r�ny�3`#C�A��l��ۚ�<�m�F|�����̰�q#U�Q���B���3����YE��+�>���YT�I����Zo���*#G��U�+`�G�L�UVh
�y����Z��g5���:������OE�V7?���qK̽��<�l
p6<gu��JQ';ɨJ7��!8E��rȰ�8:>%��E�d�e?�$�zl�����pu�A72:�Q���(��<A6)����N5y .��m�٨$����k[���N�%��k_MQK�"��Et�=;�<(�+��섶�h�������Ӹ�J§�O7E��/YE�#/��=��.?G����md!0�� #-k�L���|�t��3=�2��EȲ�����y���������gƍ�QἃY˘����Ya�^s�]��!�\�ʏ���3��s���!��ן�ZC豆�ǈ��O��,�������BGkH��n��}Э�2�qo���(ؿ&A���1.��
�HI�2k��AS~�l�*	=:>�5����l*�"�����K��������+�m���@ݴg��?�z��#99a��"S�-_
��r�1�d�fj��vaTd�6[�`,,��?��9����1ĳ&ּ��@d,d�8���Z��N(������h��׾���*��d�K:�6ʺ�h��W�H~�8����]���=�o,s8ٟa��'3�6_�r����4Ű\g��8z�3����5�E���N��1�?jz��+j�zVŜ���t�̞;_�<P6b�*�L> f��"�(��#��,Zk�6\��y}Zkr�}AQ�����zZ�9lm��B���|VG��6}�үu~\�_�h��߯����L��1_=�\p𰧄e��㏩�GmE�֏$������g�Pm��^��i��K\\�{���"3�~�%���Ե
���vy~��~�\�5�����'�,J_�Q�R"X<�{1��?�jֲ���w�/�%<S Q�|ڗ��,�����ED�blj�a
/3>�.��VNv�ѩ1�V�T"�&O���H)��/��{�W�;���a-�g�ʝwh��ɺ#6e�|K��JJ��kr_���o��8��b7L>��. ֯V6v�/���I���-��/�{��f�������D���;�%Ί�M���u�{C��r���%��Z� ��9m6/�|�޴@�j#n"�Ū�%�9b�2m�'���n�܁
ŁY�,���iF�]c9��@ɣ�d=ZF5��t��>v��R����Gm�P���h�Ӹ����|+�X��r-�Z3^�[�n�����i�"����)�e�����^sw��؄ݣ�(�)����S�J���Ր��4�cf���:�ME(���j��h��S��x��R��KoSy�J�&z�n������J��Vv�GI��/���� 4�_�}|@`�z�9h��!�0_���vY�Ѱ2l�=خ���.�Z�%ꨈ�NK9F��A�zf�6�`�(i��.'1d!K'.K�(H��OF�7�y�Ko�.���Z#WA��A�˫�(�B���9~��述3@����t���ω��68���ԅc�� g��k	ܺr[	ͻɂ\@���nu>�����u7���"��'�]7��֣��=����p�%��Yn��#���7���r�Z6�"�On��5p�ӗ/��<�3����Q)��j?֩�y�h$n8oxA{��o/�8��8��ƀ���5Ɂ��p�f6���5ܦZ��\��y��%��� 3`�_'1��*��NwI�Al�~=ifYL�
�|���Ll��z�U
NG�h�e�K���MWsŨ����V|J�ɢ���M�i��`h)GO�˷K���-P�3j�O��pJ�9�J�i��22Ԏ#�*�p��R��BR�_K������DĂutn�k��L9����Ӯ`��p
R��C�B����Rq�ϮFZ���"r�����q��9r�G�dƖ�#�f�`J�0��44e�'�.�T�M��z?�0�awC�B�ޝqٚ�.S	su�P�1�hU�l���U��b��U	�'�7�bJ�'��V���>c�0_��i���/A��#��w7˯悏�2��>_�m�B�)�-�5UN��/�0�F�}[�#�w�]�0y�ǪB����g���MB��x$��װ�ugX��(�D틊	~~�?�3(%vk^.����gĭ�Ra#aU���\��c�IM,�v�:�MdB�	��C��!Y�zfi�S�5�V͑.@s|��Ai��@�dޤ|)�P�:��B�B��985�>�`�]�>�{�{�.���Z�_k���$�,�cy�/QTGR892�ݑX5� ��������q�ך�c3���/�%��oQ�n�l��_]j�S����Ѓ6XT�{������oC�N�;O��Q����~�r)$�o/�f;;��N���1�v��Ku���(���-yS����_j�KX:�ʛ���5f�YݝaS��Ґ��������Lؼ�V �̏q��i�d�@�}NKZ(D��1�*�\�CE�v8;��[����7`�������!=f��b/0������%�x|�G��=$2$���\q�(�>�����%���Jk��c���9�Q˼����-�rʃ�_��㮑y��p!���7�皉�ϓB ���eؼ79?���j]S]yL�W��Yk�TH~���w�A7�9�����@��@Ĉ��=��{ϱ�XC[{	���{�4�C�	��ZM�� ��b?���+���D`��LuV�}� ŋ+�D����K�s��uN����;S�D��R�Q�/�}��BW*��R�[�Ǜ=�N���g!N�3�zg~X7��F���_^�9���U}a�I~���(�	�rX��"��6�|������Ta�ey�%Q���6k���焄B@.u\��0�I�"���N��a�Ee�:T������k�(�II1�b�����e��
�@=����s��c��*���~��?Y�[�8���Eg��`�b���3���ky"�HО�Ա��V�C���ǭ~|<4�k���@7�]b�ƫ�X�D{����SEF\����hlcq�r�6��큱;0�>��`�]� "�3Otf��=6�O���"�視O�ŊV���%���<�*���F�5�:�QP�MI�r����@���0�"!�fhGR�8t�꭭M��Nx���8}�h�N@�Y�d�w�l�l1�]#o���4�,px�M�b��cg���i�����0�
�-��'�w�� {u ��<��y_%�1<ʐ��㠶��fx[]n;
��L��F���5Qt$	��L?.p�;'t�^�@���)v��U���LF��`�=2�TEZ�F��E��+'"��2��@u]WH�Cx�x�?O�́��'�&�xyv�
�NO�k1��"����n��������.�r/Rd:Î6���u��©Flр:�wѐ�;��x�ɯغ�ģ��Vc�s.ac�~(!��+�����[�	�wW��&���?�|����]�7����m��Fk��D����K��\�FZ!�*?�H����2:x�#F�H0��S������em��(�㼦3�ӉF���Kjֵ��nƉ�=Il�!��d���y����~��sT��*�����}�H��Q�'Q�:�ė���f��U0(D.X��̵f��K{ia ��a�.%\��ihsW6|FR�(��B��D��8R@��&��6�C�:��އ�>���gp����Æ ��@�z�/4V��RD�ك�Z 7���M�{�hW�� Z�L]}�ƥ�<U��Y��E)5�a��\�~8�8	�<7���(�;a�(-t�I�C�P����+X�a��̒�b.<L@p�X�����������5�	�$�x�q�>��DJ��~NIJQ%�i���.��cF����}��Nt��u�^��R�����FC}�+������7)�ӹ��`�!��n�Pv�L[��@D^����n_��ϼV��/�L/4<:��-�d>�>��2v�g���b_���sD�}��ɗ����z�A Z���F6`<�}�yGdk���P`=�+V�Gk[�^�eN��_V��n��^�>
�
2�7-�r��l��PqzW#\�C/	��֟�ڙ���rJ.
�S4�gß���d �l�g�;ύK�}����P�&C!��h%�ߒ�{����)Gt۽��Ub�\�3��&'�l���-T�P e6䲎�Q�P���Ya~�b๏����YТ ؕ��}���եϣˤ}f��0a�ftM������h����m�k0�d����X�C)�^�〕�d�Yc�;,�D��Q�o�1�ˎy�;r��6�z��!�e�)�g���Jm�����-zxY��`����"f���P��f�A8ĜF>BiJ���b'؈=�{pNj��V�"ڱ*xH3����âDUk�(7��@�35���!���κ5�+[��T�W���k�¥�mJ!��+y��A��J�C�7e��$�t�js�E�	��" D���9H�j��nn�:��Gxk�Ή �k �h|���Y�Tc	7��~�ʕc�]m S��5{I%�܅�A	���y@0�UR>�F�R��F2���H#�*P���W�Ķ8E^n[ӊ́��$�S$;T�
�cQ��q�0�����(��q�Z$���� ��hQ�<�ݲ;���zJqپ�%Tξ���'����iv�t;j�v���?�{eġ(�%Me|74W}��{�|�4����2Q
A�*n4)q򝠷�?��h�/�2j��r��C��x�j��#G��f�$ ����+��W�i�T��y
#�:4��\n�q�ژa;�t�vF-
��#s����[j�����G,�kf�灤V�p�XlxV64EB    a1f8    1b70�7�A�|����R��w�e���Ƀv�5���-���l��5��W��y�8��0_���O��e&�*��u��R�Q�"��"vHQ��nKk]Î���R�F�+,]��[�r$Y�;�*B2d=Ж�Pd�����N�����/sQ��3�@�K��(P$5�0�9��-����Cd����D����o��K�4�A������1��<h�3s��Ψ�����h�j7Ͱ3TX��Fx-(zy�� �����$Լ�9-�-����T@��#�x�H%%wc�ͫ�B7y����1�hPQ�f�<D�WΦB�!�����ߗح܂�at������,Ɉƹť���i���AnUv��Px�'���f�tðd���ّ�˵�at�[��gMɅU��JɊ��N��׸u
~z9��ޜ-���\I~ζ�E7ts���j�-hX�逨�|]�y� ��l+�O᝝��o~�xkf��S�Q��Ƈ�N��.���xñ��<�R�yu1���T7M{����P�R��`����?M��^3��|H�`�܌������R(9pW�r���1�OqP)(| �y3���SCz~�K�oQ�Q�I�|N}2w�3�B)���-�{�W�������̉��%�D�L}��ȭ^��e���PR`��x�6N�>Thu��N��� �U�W��RD^*r�<2z�������tzxY���#m��  �0j摾�Gǫ��@<#��O�&�ߒ�J�Ҿ �-�O���B�]���D����\bU��ц���)]��$h�����:�������Ba]���53�i2Me���h�S����y+$@��T.�M<I8�6=m��^����;����"h#�|��sG��w"����D���3�W��004S���񚓊P�,}u�;qn����P9D�l��o����w�Ȭ�ŏƬ�5�'ʡ�>�6�7�o�^��y�aH4oTu��G����(^~]D�g^�r-3{Ď~��ζ��� eE��w6t';�w�Lf�L�2eR.���+���k����}u�� �����@"`�r�`�y'�I�&�����I�*y�o�,:A�heXΖ�l
n�i�NO*�祖��qE�n����*���,��N�UhG+"q	(Ȑ�W�o�P��D�=Щ���1w�����_���G
�C�`MX�FJ킿WKYdio�������ܝ�"�[E����
�Q08�.87g@e�<56�4*7M��t#SC����Y'�~���Imoc��s�z,g����ٿ�:�@9 ��O���8��c��W�,�K#�!n�u��Wj���fs�Y���x�:�H[�Q�S|B2��WU���?EBK�G����� �x�Ҧ߈>�m�Y�(�>���f�B3p_���h�*����Z���@��8�7,]<�+��w��E�-[�KL˱[xUf&7+W�dRxFRQ˧�IM�8ݫ8w�h��{^�vFU*r')���o<!A��
�)��OG_�����n궎A�y�V0�:%�G2?�����݀���{�,��*J:�0�Ixr���F��x,1	H�Jj�W�������q�;)����qu�Y��F��Ff�fQ)�����U � ;�C������v���#��'H������os��"��6����tB�v܅�
2�Ue�h�KI�jG�_wE���$Q�� �Ѹ��(����0����Y�Y�w����F�?��ݻ��-ع��Y��N��J�O�f��_��I�.���7��U0G��ru�o��F�Xf�a��Z�X�[#?�Y�xϡA� cO�1��G��d��ߙ��ݾ�!e�0�J/�h�w5�����B�����fy�=}��	37}\�~~t3c*8m͎X�kn֜�;�eI�RN�:ǲõ,�]ү9���<n�+�|m���V|\,فA؆p���#琴�L0t����O����s["(ed-F�p�ꃫ6�����6�kĨ���H�\˰1�;��=����	�s�gv���3���)d�4��`����A � p�֐G�7�D���-�>"��2[U��FÈ'ɝ'E���y��=�yqI���C�嚏���������o�}���s.�{�uMl��2��K�PQZXR���ĕGޕ����P@�|��(_��3���Hc�R׳W�c�2$�ô��Õ!�$.�G��dú�^Db�ϝ'j��3���VKm�.;�26lY��,�8P��N�n��:�"$f���a��]��o:���n(˯H�f��4�N8�\ʿz�1�����`��`@d��X|���=�f�e._�����ƫ͞���;lNR���!֒O#R:.����Me���vP�T^�~@�]��e�N��z"��}(@��&�����`�Xc���=[��@C��o��=��ӰA6MS�:����Դ��^
G��a	ZB�`<�	$:A�a�%]��/�Iٮ�R/KGs_xd��3Ѕy4��l'��UR�tE!y[�i�"�-k��F�_P���/H�h[��`z��)4�K���o�C�����������(�(j$��r�ʩ׸DZ���i|B�w��1bq��_~N�������X�nbF��+�}E|b��=+!\;��*�.uI��kn�P���ut��i0o���hd��O�Z&"��W�21~�.�nx5����(D��'����9Y��<j�L�Q0�F|]���p�ѥT"�Em{��5�r�����R$�i�����)V��^�),����*�t�~��j�YǿkZ.�ĸ��>����
��;U �Խ�H$xh�'���0
QUγ�� �D��S��_��M ��ٝ���@�V���Ԥ���݊��G�x\��n��5����d�H4�>c�.����N?��MH�pMv�p����r)PK��k%��xBdB����{5i��|�!��)u�K�t.��&�*��''����x� ��z搥Z�8 ��˼j���{���[�t3�т�LVIͰ���-2�j���aT"l�+ɷ���I�ڣ$J��:)�����v���h(A���ڏ�������e���0��t��nR����� Ø� �|�.t}r�������8������d����c�vk�߭�_�8���цvoM�\��!�:�jO�����/)	<;W=�<5
2�yP_���sm�[%��fi�^�HohBn�����?��nt��w'g�2y}	�I��8�Wb��u�U��J/R!|�d;���{v,�@�?�Ӊ%�q髫�E��U���+/I����`�Fũ�gO�D��9�
u�BӒ��0�j�b�a�"���OzW�<�`:���(Η��Q�l����.M2c�O��n�l�Z���փ��1m����@0m���6�p 2�TDC;H�-�)�>5�S	v��)�!d����|7��x4"R��XY��<����<𬞣�H������ chU���
�)-���P�2�x�	�o�̧����Ͼ���"�V+��[�(gU��"ƻ�>C2�sﾨ�FVӴYq_&�L�����f��8��*"uˀ�����ϡ��C��>�~C}=r�(���~�O�[�"c���:V��y�VN�}sHyC�?��_È�A8T+%�(�v	yn������>�(�`3����vDMfݲ�ɖ�����W��7���e�����µl=8�$³��U�Cg~�Z�,
dnc�( ,��:�?�c��a�c%0	��\ #�x�"^p���|����RFO��W��Q���f�JA�rF�kD,�C˵����XR��C���r����$�Yrۏd��"$�u3A
lyސ�U�Sկ��9f���o�����f3�s<CD l�`����eCA�M˦ފ!wo�x+B}XB�+�i2��0@.�e�
����D�l��8��_�	�l���(\fO�iwC[���J{]�u�$�ݗ�}�^�V�ڍ����T���h*�|.�c������S񚑀��,�3M�k(�y#
z�=.I4UN�(��|tH�&I-OQZ0�0��K:v�',-tHM!w{vݖ��)[y�������3&���[4`K��1$ё���#��1�;`�C��́���G��ح��4�f���C�+Z�\;��>]�hP�?��Yd�9k�
$j���Z鷄.ç\w�3���)���]��%��8�*��_�|���H�����v�K��C�����3Ə�>�0\g�e���(L�Ed�6SX����%�PYK�/�N��\��$�zeQ2�A6�e�+t�n�H�ݻ�װs=`s'9�qY����������r�¦����l$ƉK��wp���-�Iʻ��~��%���d��(��ՄO����<ۯ�ZG�^gH��n!-R�-�8d�!���#���ں5c�5I��$���(88sg?�`Z�~�iV��k�������`$T��[�n?�mq%����˙ȁ�ka��C���T��!��:�{��V�0�&�sĒ�=����?J;�w�j7He�����g���[�'BYe���Vmj�$�i	g0e0��S7M5���e��4�V�� �̊��Þ��c�+ �mɽ��D��L�Q%��}��`�ü=O	L��-��P	��vW��陽�g�V�brJ�TqV�O�f	-eϬ����T��L}�Ԉ�1�/E;�ү�v�������(y�������ۇ}iY�}�|� Y�8�wœ��?�v��Z����5�ƥ-�'a�07��6H�>������S��zt�;FT���Щ�;旆���-�JH,m��IH�ٰ�Ɩ�_��4����ˈ�b�����h�k<g���H<O����W~��9v C�\���n��G��+���3v��?W\cE��0B�_�>��Q��X��?~�XK������Ps��H�(n�'�a����rڪأWv���;Qk%�dI���A�/�gO^�j�1� �J5�1�`���8̳][At�L�]�j���_[S9�M�)c���uv��1�9V^�
�;�*11Uј^h&�(�����Rgi�05�A�/�5IJiw�[כ�r�[�K��F-����+m��\�Y��up
�l��B��%
���a�1�T�� hd�cB���	�)k�_~TL�=���s��6[���Y��-�Q��r�ґ��R9^N@�4G�
Q[��k֐b��Q���D[>2 �+�	,-�~P��1Y놮/���p�����7��X��Y���F�#�|��P������G)k[ڞ̷�z�Ȉ��A>Uҍ6��m��]��I��l�\��w~����QW����0w`��s��7�(��.i���m�e��H��[8�1�;�"���
%��б2|��#/=:�bz�Å>�]��F����7�c�;�&?�������0
ʭi��_�!m��g�]�uu�D��������I���vI�ŔTq��w锗Ꮊ"D=�ٚ[�l�J��Q���t�>�����*�32+s���>t�Ї�W �~�>����zS�g1$S�	z�4���I �i����y�
��(��6*Xb}�Iɕ����M��X��xY��S�m���u'��ң̌��«x�O�5l{]���> o�^^�ax�	���sYÌ����e;�=������Y�Y�W����
�K�/�����U�a�\E�dL@��u����ȡ<#>L�V$��O��OuYH:��w���"|9K9��8AF�k�0�=^�U����n`�B��,�k�1i?vF�,�H�]I�K�L�/X?�2�a��}H��m���V6ź�q��3������:2���Z����&���U�TЅ�Ư*�������F��D�_o�P�Y���Č���R�������F��o>�0x)m`���i��������%_�ſ^j�}�ҧױ�g탴���p~�/��mF�ȕ%@�]�o�/��V��](3N�Yk�}�?j�v��0�:�捜}�7u�������ڼ9��㢫�c����H��Ն�I�,Wi�w?]$�w�B%�������샴��?&�I�{C����Y8��<hQ���å&�[�[á����J5�m�Jt��x+r������HZh�����nemd��E�V������r�����  hrF�ƨ��� gE���.�:��똒���PS{�u} E�J�d(�����yL�ޏ�ztvjq8���Do��l3�Z,��m���
4V�"�kNb\aG�B#>#.ׁ)-�1X�_AƷ����G�S��x;G/F��o�?A4|�<8��G��4V(m�ۏ���>y�VyFM�{tb���d��t<r�g�`�1WMZi��[����̕w��gf�bxF�Y���|J0��pN���l��&���U�Q)�~��l(�(�S�Z���Q[�áu(��G�~B"�$���|F��Ɓ�q�)�H��%ಀ\��g�g鼸����S���1���D�D�ƞZ�S����^8�^	�q3 |$�Cc�Ϝ=�M���n�%�m3y����q��	�=u�]͊�zΎ���2RW�g�~}~!�D��O��O�1��UH*�b����s:�Y��`F���y&>�c:[��k.(�S>�Ǖ?)�#G�@�\[3tԸ�ЫI^tJ��T3s,@��y�)=�!����^�3%�1U�9�Gx���$b�aG~ºd-��$c�Rt�����є5�5�CR���������ܔ��,���$U�e�ea$���o��!�$�<^Ǥ�]6Ht�@���W��4�.� ��6����]�����H�.6�����_���!Ru"0��E ?C���r�]��5㶠QJ���� ��c*?�.5>�.�� �Q����)�K�2Ҝ�����߿��p�I�J��C����S|�,��]�cu�2�*D�C�)i�wl�@<�ÛY��6��V�`���D"�c M5�