XlxV64EB    15bf     850Ό�O��K�X.�Մq�>j^E�����_��sװ�=J \)�F,4,�b��g5�N~�T)��������.��v���p��B��Kl$1�0�-�G߲T�Q}�#�*1�o�u��V<�������eW��N�Zې�ci-�3bs}�f���ʻ%�v��K��o'i��M��1�/#�?r�G��ޡx>󐷈��w]،;�.n@k�'$"�D$av�q?�)>�E�� T��D�h�]�?F6oS,�}�%��O���Tl���y�7)gސb
���)���"���S��V�
@�:��]	l�)(����1����"Yɭ���&ih��Ő� &�Y�+���٤Zl��4�[�-�-F{�X�����AO����]�Yۢ�?d���7E|�,�������= �yL�X�n}%ߧ����c�'��o��ZnR-����x -�G�!.�R�V$���u݁�s v�C�ģ�QWq���L☵��>27���s~�-+-��U�������B���}K�'C� b�S���ʖY�ox�;�(؉qJN�'w�@P�>�<��
�7�V~���:b`Ь ϭ@U<\r�)��X�:Z���oYfOu�9��ڐ�P�6�*�Z/��� �09�Ȑ���u�%����ݏ	M�iC��ew���~Ťl��!��7���^8u�� ݈R�\/e7A[�hZ�����Vo³gCd("�C�XD�D�,	�"��U;��"���~4���ΈW�,W���;��0Z�p�eg�<(��E��^Y
T2��������#�B�\N)��l�
�ɂ%�@�JĠI�C��F?�m��R��/`��P�Lx�%h� ��$��7��5���~�V�~���JI�h�_��#��菜�=3�����=
�8j�?w1!�W<=쀄���0 �Y�t��x�:p�ko;�8�+-��P��XsU&�������5֝m�Qk�&�X�&ЗJٕ�Hh�J�_�!omsF�<�ie����+�U$쒢������*���ؿ�.��$�湯`��]8'����#s�Ж(�Q��h]��P��N�_�0c�O^[�64%}ao�l-N,0�<��,WluG�3��U��<OB��}��M��d��6ԍM��j!]�o�W ��+���c�}$�� pͰPP0�T���͗���������������K��Y�TO#�n��ێ
�n���g�gs��Q��k�U�O)������߭�z߉��!�=�?�e���J�����`D�0|P��È;�7��T#`��r�K��c����Z��1H�1��H4D~+��� f�\�!��|�:�m���z�����bqxI��Ģ�n�:����{8箛���bRT��8Hz����T��b))��e��($�,6M����;8~�.t?��~��eyVg�]Ĝ;�7��b��i	s�`,))0����;珼sֲ� �7~8&1[��}je�ɉ���J �O�K�G��X� �W�̶�z�~�f�&�q;Ϛ=�F��Jٓ�[>-^����a�"�9�|�y9��r<�/1o��N���u���i *����Q�/w��Uć�6�C��;m�G?\�Yq�'��[� ��n�Ҹo0a,�g��l;UZ�[�i��(%���VDc��.1$߁��q"�/x���+������(�J딂��?L�{�� ;��⯔�O��������fZ
�S}��a��;̜��y����&Ru��F��q	g\D!����d��+}��=�^Mդn!�F�Ky�<�o7踒�[�W��&J�#���Y"�
�hM��WIf�� �_��;Jt��Tmk�N�q³N�^U<��@���]�O����u�+8���9�+�AUwB7�G�	 C����_n�f5��O���)|����qȾ�������!?���55׸b:P��zS�!��0�13:�ZNY��\P��|�O�2^��'ݳ�s轹k�ae"�(��z�O��Xǯ���;�ć�f��W|��Ό�n�_
�n%��~]��pv����oH�2c�S�Æ]�H����pC�V���=|�E��`���y]�Ĝ�0z�21��>Z?L\�S��U=�r���