XlxV64EB    fa00    22f0��\,>��kk�C�ZX�5J��5��'�7.��m���*�Т��FPd�7�Į����*[J�k��SE[��v��W
�RX�%�p�(ڸ4<�y�=�8�RN3��S^~/��(��*��>�R<ؗj̡U�%��C�{�����7U$;��#��x�8����R��WϽ$w�d1 �V	閈��?މ=��9��T(oݰ�4"�Ce��4nK�0('x���J]�Q$\K[�!]�*��j��>�� &WE�]3��s��'FU�Z9��6e4P���~���ó���V B�%����{��%�Pz� ��L߇��j_eLOG�,�3��{��Ö$5��*��X��7�a�Tk���S�ӵ�fth%�eQ����[�C�л�Θ��� �?-�lD���J5�idPPx3.�V��cg\�����X*��*@�ʩ'.�����L��G����'�����S�ӈ6��B @�_���[��x����`VM�$�q���:9�-���='0.h��b1ы��^4E#$�>�rЖ16��:��-/�|������~-p�]���j\/�_M�'S�T�c!�Om�]��=l���a_�\ws�&��N%�<��-��܇w�z)W�*F='V�5�����L�3qǡ7?jmp�T�v�����p:�W-U��&Io2�8��8������4̈����^RzaZ>R�
����}�P���ْ|Mg�5�e���7!�3�7����ގ:�|�mn��ma��!�01�̓;4����A���?!�n�@F��\HA1+:��4�}Zt�]���I�ǐ����Z!y�j�߹���!�'=!IV����[H��i����^c��Hc����$�\���ǻ��ѹ���6{p��	�W(�!���o��bD�]j�h�J旸L$zwm:�n1���tؓ<��0S* fg#�nvh��u�&�PXO�^)�R����������N��)h���N��{9�-#�*7K�"��(�p��"R���.UEB"� Rp�h��u����'����b\q��R{�~��M����)m���	=�+;*M�s��=�slkG�B����>b4��J¨C�
�`<J:�ǒW���
���f�^4��m`� �H�|�����5�7�~Ʃ���{�.x��C�L�q�m�6�7)�ۡǽ�5��s#\��j�<�%i��5K��v��^�E�C� ��X�.�X` �Ծsp[�QA���&Wl����/~����s>���Y��8�CQd5���?�9!0��OR���ȯ�gW�0�:�:��~7�N-�6� ��	~��N��,ShQ���u��r��N��h�*<��H���Fo�H�(p'��}��
 ��b"�Sy�Y̓��[���	D�a�aW{�t="*<�)m��Ρ�~[�F�o�̓��m��*Mv�Ȩ���A����0�m��̠��/�9�&!i�e����d��C.�I�:�H3��ȋ� D0s�.��=c�!CME=զ���53nX�"��.z�<e+䫮�\+��A��u�����EM"w���-�'�ėZ��x��±;�d�]������v�m�U{L��F��N����7�%��;h����,x*�E�ُ�Xı�ҷ��n79���N�e-F��f�,TC��_E�P��s��7�ћO�)R��L��� ����u�!cC�/2�Q�V\���)�ɾ���e�܊6�l�3}�H |(�҆�W�����*�L�r�'�� \��jJ<�����@�m��!���������pMè
���u���A0�qP^�z�huS��p"�G�k@�@X���K�d�Kl	hQwXPL��X����O`�����]�V�ëva���<WbCc�>�f�	� �-�"N��[��a9q����yWh~k��bu��yu2��8��*�Ƨ���3�]-ʹ����P$�Yp�Ʌ�!�Ah���b�st
����[�h�Í�!�gp������,s��eF���.���UG�~$��Ј�}}�&�]��Ǳ]��.�N�~���-��8��p�D�b�@�iF�ۉ �sP����%7��s���6�L���VOA��3F���`�+���cɞe]��!a^e�*w�v�F|�e�ʝ���"�Kg=��))B�?�ɧ'�B�gͨe���9x�姏P�l����kľ�l���h���� ��!j�T�Xhj��::A���`�^��OFR�4<��bi���l���r��7C�� �ȳ���G�F��Pּ��I˷%�ߋi}��t��K��5r7������ٲ\�IȆ�	w���}30�Rj�97�����OC�{�J�.J�\�aW�F4���i'"e�Y��J�G���
��P#�#Wm��Q�F�KZgU�MɈeo=V���0p+B�R|��"oRH�u�㷳�y�Gɺg�U��\�
WŽ��݀�:[��u��^���kӫc��p����~�/!���%`WbY��_����tp'��&e`X����z�����u�h7-��e�.�\C�U�(3�����z>�I�S�-�>�� ,�rpY�m.����t;'&	�$�����#����bm1؛��	�S��0�Syl:����i	ҡ��ma��r�����Uo�)kI�]D_y���ܒ@���$��i禊�F��6<��c����рR �L�eƷ:����o8jB�C�~��I��Oʨ2酨jINNvu��dq1�3����3�Ӣ�d����F�_�T[{x@��ϔ]�4�#�����_v]6UA��n�I@��� �ks���Kx��k�R$^Z>9�q�>��`���q�KVF�;��NH�� ]�J�9����s��-�]^�_�_y�V3����^ @ӕ��P8�ے���G��n?����P�N'��mL����� F͍�@�B���sY�^ɫ&�Ī��=e�7p��Hxx�Յp��"��J����^��vj?�������s��DD�: �R�\+�r�kq��z�DG��Vp$�<��u���`$��sK�A����	�9w��w�^�~��4�`#I=��d���#�mO&*����*u��DDEx(�5z�:QO����X,-���.��iǋ�my
�`�YY4���,����*m�]d�������Df
f���C? <#Q]���B���x�i��BW���ա�Ʒ���$e��� ��3xy�s�"�H�H�=O_3bG'�j�!�e'�ZP]�<VO��d�/
������>Q�u���iO��oֶ�%�k�L�^�20��]��GNA��8���ȕ���O�A��O�wM������O��������U5�^fܶ��ع �e��3^rh:��D�ß�sȉ#�v%�T�A�'�7��0@��r
�yH�����1>�;��������ۯ��fb�t�T|�	��x�Ӝ������5�M^{�����_��p�·J��is�(�"�� Q$>BB~:���L��ev��䧑�:�nHg<�fՁ$}~����~>j��3/�����7IӺ�NI%���kR�����) ?|'��v��o@��uy>}���d>^��E�(;eU�ǸU� �)��K,A}�u�����6�&�(���ߤ5��0>���,��pe,��M�j�[��n���-��w�����d����p�:�{���?���STZOJ��J
��X�Ğ� ��r%@R_��>�x�~8b4-�V������3�4oe9Ae؎Z�68��_p���I쏡��{/w��b��:q$�ͽ]@tEw��c���X������T��*����2E���k�*fE�y��O,����+G�3x��H�\N�>�h�i�VkK1h�H��!�	ӄa?�ے�C濮~r�b¨lNA"-54qk2�����Ʃ�s��:�m�GL���Z^���	B �	J!�F�o�
�F�V�����]�qk�k@���X�h3��P>���ڜa���W�`}�uVl�s�\Gw��hE�W��Ybm���2I�C�[��x���}` �I�����9e]�K��|��K;��C�$���?�b	���E�x�Z�=�iV*>X:�j��������X�qd�i]���e\d �yW�{,�=6򸲲���D�?�|oM�ʵ� �x�c~�,�A��Oe$�z�%��������[���eC�x�����~�|=6,�x���񐞳u�3�H�ͫ�ҬOQ�ʡB�7���N�M=�}�|��K�Zy���,�9����A˒�-&.I��P���Z!�D�:N�����hK)m�+i����4`L�{EchϠ����Җ���x07wB��cp�L�h�^Nwjd�{�4dWv�^�;�E�yKކ�{ՙc��R7�wy@uHׇ�/�8�x�VBx�tʿ�\M�Q�њ�~3�B���bLZ&�/X��)�-��	��@�ޮ=8�*Q��:"�利sQ�<0�<C/柔�-�M;�y�_��A������(N���fF��"���=
��{m��D��)'e*�4X�;sŪ>"��D��� 
%7�;�7]B#������{5��Jϊ^�Q��"��~ݮ�/�6a(�CS�1�����DD�>�2��pG;�D���o� ��m�v�Fc7���YL�_�װe�2��A��Z,�����#��=BqeKϪ]! ���{*2iX��lXZ(���x�c-�:sEqu��E�\I:�!���扜
�0��l,Μ��K�9��9��C�@5W��<"ӅW��_���k��_�&����V`���.|d�H4�#f�������M��=U��R"��7�F$�pM�M G�I�s�1�����Z���4~�i��D{�;ޒ|�j{�U���˞+�,����Oj����d
Tw.�הj]&�'-5��x�J���#��pJ�gC��f�02���:�z6���~(�-��GT�5<&֞Y�9y�R�"5R����g"--�"@ި׌�s��;��qb8�~2B'�sxT &U��!���t�T~@d����?QN�)G�j�H=����iS��4�}�M^����*���
���>%�~��m��F�Fe��������?+>��v(��������lLS�����GX�1ki�Y9Z��yO��pz����3�d���l�B7~�5�X���bN<	��h�(o�_��~y�"n�\}*�!�&��q��H��J+r���:4���� �������>����_�n�a��Rkv8a���/���4�.�c��L�ݵ�gJ���M��MObm��1u��І�J*F�nZ�UD�h�<GM�NP;{��=_�}����Y�\�Y��#ly��T��ZK�Nb>`K]@��i9�>C��c:.���_��9<el��`��:zJ�l�c�w��wu����:cHp����=Tj�J*�wZ�P�ɠ<=ˁ�����w��+��(�VX���MUk�0w�%�:�K��:�R��	x����C��M��{Z躉�����DKf�D�[����hm_[{�Qݠq�N;����8���o�ʇ��&D��T�yB?P^��^�N�� C������+}7��YJ=>�b�T���A]���f��=��7t����ǽn�2߅����bYk�V��c_�/]���!���O��0�1ʠxN�/�*�|��߲n=�����}�
�T� ��ԨL�2�g����6�w�og�Xǔ�O�ܚ�1�m�@�E��P��#�:u%��Fp�.���"~3�� ���G�@GĢG �S�����n�<�.P��M��P_���@�W���}��^ю�X.��ag�¬�����Xaо|�^�E���iY����P�Ҫ,����Q�x�`�����2͉H@Ȼ����CtJ�nTgu�Иn+����/���U���jT����<�zZ����-ƽ/��c\/��{9#�������E�!��|�}����:@w�P_�qC��f���b^�8��Ͽ�bI[�rp�o9�`�c��u���|
��|΍��>�Z��*O"���H���2�Q� A�J�R����8��ѭD�و������m��H��T���Z�^Tu�)�Κ@�{��ZdoF���΁#�90�I=V;��&�Y����5���9�yT�Ϣ`�__���BI �����!U�弗�>�'�u^���O���%�o]Ղ�{LJg�;qu+���;�&�-��ޔ�waf�����jE�����}KZo�]�*���Ѓ"av���>q^�x�{���v��LOOge]p�B^��t��=9-)u^��ޝ` /��8n�����e1�YΪ� É%��V2I�����h��A�K��5���)����-�L�^c�f�{�E)Uk�)g�͘�p��i������ �����f��R~s��91������!G�ʡ��<����%��h���	�+d�S�(��p�v�^<�bR�BJ_(���J8�O(��KI�Ax���q�r�>�0�����o��0J�f��o�_@�~o��32Y�<v�R����9Fiؕ6�|'�ܫP���(읇	�X��+WX#}JRD1/��{B�ɉ�Ρ
��6�ℿ�$Dz�c�ihgdt�~���uP�Z����~�/��S>a2O�b4�����k�A2�R�S	ŭ�fy�7���99oL�5�ܧ����I�St�x��zǛuiW����AIX7�2LW��(E {U�B����3z�Mj���� ��9z��q�Z�Z��X����ݼ��%�
׋ ��2|�9
?�������*Y�R����a�C1�Em����(K��4:d��4<d��G$�}/���;g�h��������I�|���V�-k`+��v�~��N��+{�İ�@��Е���K�����h"칽R�>��'��l��� ��o�|H��9ȝ?�^.j|���V��vYB�/�>
�k\��>&	Ac6;�"��U��FSi@�#�K�ND`�H�Tj:�6�J�/C��o���/�� �p�%ٛ���GG0�����L��2Mx!�{�����n�iW����D�`6�*]1t��8�7B���}w�f��Y���������z���CXT�<�M~H�0������0�m8�(������XL�Ϸ�J=���˰�+���V4š���.&�B:��D^&O�^�9ZKcd�'dO�f����\
?$Mb4�0�6����<���N��S�VmZ[jNٟ�ٯ�Ħ���0�* ��a�≯���g��o;dg���+���V9��p��&3�BDd���9��2�[��H�2x������7�Z�3�Ô�\4'��>��<YOi��[oI���w�-}��;����>?��B�c�+&���C&p%��7?� ���������i<�j�:w��m^&M�]�>����6�z�/L�'y���͂�-�!��#�h��C��Z���+P��{�#��/���?�t�W/�3�^����0�U��dO�H�Kf�`G#�����>/z5tx`4K5K��Gg)��4߁�`&;����I[u�ζ?n3�T� ��tfƪ>�T�\B� ��C=�yq�
J�}8�]r��:��Gx�G/�v����2Th_W�̑QB�n.Jg��S�}1��T]յ\�o�qﮛr��cl��
#̖�?���{�����6������e_����U��.�Z�H`hڭX���G-������Ǚ�s�e��*`zDZA�Ȼߜ�fӎ�]\��A%΁��{a|��	P�O�h8�k�zPs��*8)<�5�<�=�D�5��Z9����9���K�J
�R�V�h�hI��N�IfP��<����%VDc7���C�'�{`,lw�o�%��O�Q��̖�2'�׃<��٠%��q�{^�� �/������\4:��8��@���I@����A>ڮGc�v�0^L!��������Ԛ4V��g��=�U�з�ͫ̂�a��� ћk�B�MmUM��f��^�*���v({�8�����2s`Я���!�<G�b�jAduy<u���(�*h_WZ�!����-���,*���(k�
����_'	�z���d9�Pj+�r�5�o�����Rc��ByXc��$�������ro0/J��dJ���^����ڏ[޿@�Mi��D
�M[���d�ɐyo�fb��W���n!��U_���Yp���%3/{�UrL�=2�k߭���)-,����Q�}�����0�ɥG��>B�md��pp ]('�7Z�/���k��^���"G��&���*�VdA]���m��p�j	��)ٺ��W���v��`��N�8�˺K���:5�4-����r�1{�e�5�t8����)�֍n���?փ,�)�)��_l���@
{涓Y�`%�n���4�һ�� Y�m���T�6�F�����D+�B���^1��4>)^;�>�������j9g?�-8e�ݻ8��RG�;�7̲���2D�����$h�i��5�`����]�Ed3蒳ژ%q�V�������'!z%a
��-P'�s��j�b¯<֖�I��!�@9�N��T;��u�� 0���2��
Z8�DO��ɪG@�v���*��P/)�U%��O�O����J�Vz*�������a��T��犺�+��&��M!ITl6-�i0\#ZU״`���i�,���d�I~5f> y�����1������a�*a{q�ʴ�L�⠜历QZ͇� [�Bš�� �0��9I�Rrx�\�a��|�ÀP��N��E�B`��H�M��#
��XlxV64EB    fa00    16e01Q�*); O#�(��"ݐ���V��<5�<Om!��놷��~5^�
�Ƽ�Q����j�`1��ƅ�69m-�I�*&���eѻ����7�@�9��G5�U�����Y	gܐ����/G�ȋM�qS�ہ`J%h
�pv���.��|�CS��gvB��÷n�
�x�U�T򥲠��u���)�+�A�*���Q߫^�pS��{�������� 扲�az��JR����t�V�U��cW3/۔�����.�_��=�����W�E��2����<1����/�๵�l��f?����Z��82��u ��z��I(L������IdE�m�XP���ޚ�t�#mS��s~�sJ��DT�<o�7$*�����Nh�sE�b_uD�Az�8Q����}�����,�����w���U�?-Tg{��>~B���[�������i��fI;<�o(-2E�L
�)$�l{G+{�-����*:|�~�Y"�tKWP{	tј�/z&U��2@�ba!l���atY;s]*J��g-�$����G��+�w��%'�B�f����r�V�cB  1@-FTAԬ�	��k7�>�lT�z�ظ�`�s�∷.�G�W�����/�����ymX�����i�f���i�h-43�����/�}�L�t��ĖZ =��|�JD���:32�MvJ��6����A�m�=&�]U����N�׮fz�v�i;�L��&ϗY��d�6�G_���`���|�Nh�9��]`���`V�X''Z�}��U\��'�2b<�E��u|B}U�륆>
{;���^:&L���_yZa�O5D�^�A�x��/7���}�����(�ZQ�?&HP_�I��������ZG�-��­�Y�eW�NR�+\�o�.�j�s(@y��8��sE�[��\���%�\�o�����A�{GR{Ή�p	���f�v���(�����]�d-���/��	T�.���?@�\5��h�M]�1 `-�\�e�>��d
Ga�}�f{
p�^$�:[��$y����j��'W�ޠ|ah(�hl&����!�m�S�6ڇub%�fC���-7>�S`�w������6#g~7���3��h崼��
$T��q�I)����O9~6-Tƥ>��Jk�T�rK:��(�\�������c?stԯ�ؤ���t"�k:a�㷁�����z���{t�*:��$)��x�0O��5Sk�
��U��W\@��8��	F�Ifm5TN���ϒ���N�5/�@$����%F��wjɇ��[I�rۋ�PҴ`�֩ǜƺ`b�4z#��T்�.�˂�V9U�z�M7g�_k9Ya�K�\��B� d:�����|�@�N)��xCѲ�r��NZ�%�ڒ�G�nvT@z�'���1�N4��KeO��v��Q�F��o�%����%�I^�>�T�&�2���Ą��L$����!�
3�Jd�K/*�Z�W%N�Q�듶�3z�3A�S�9@��(����J(;X��ȑ��4�+8��:Y�m��h��X�W�#�w%=
����_a�k Hn�^�wcQ�i�?HO��N��@��ľo0�u�pZ�
���.�7@UW�i�ϭ^����?��ۋ�i �: ��V�vf��q��5S��Tx�J����]�;�̞=ב��7���Q�btU� ��j���-�hHn������F���3$�SZ�`e� �R�J>�t���Е�rb��,$�� �0�鹡&u�\�'���6�S5O�ޯ�ع���0׵9�Ɯ�7��]��D4�ڋ�����]@��HG9��k.�$�<޳�S�[��E��r{������k�gU@����j8���Q�yT\�SI���fx����¯��5W7���n��p�Uz���
x��g�Z�W*n]��=�6ݵ�=N3)~�C��Lb�۪�܅3k�'!��T/�*3�,�+[#�2C��eb]��R�u��ɵ�v���,�J&���1Y����O�֖�0`j�!�	�
�7���B��Y�X����+:ow��Qۮp�/<�fq������<[�n���[�%o�Z�%�i+(�0fi�R�I'"	�7�f��*Y�C��P �9��<��<�đX��כ��DM`��Ԏ�&�3�q�ܲC)rn�R�~ۭ��4d�N%(�r]rq��+p��5p����{���D���K[$���o�HQ&��z�,�{��wY �:B�sz�(x����J���R��z�ؚpɖ[�E�ʫ�SwĊ��e�.�3�m}��M-��ʰM©hrn�d�<�_�Ŋ�Uw+w^�5��X�?�� �����pH�s��v�[�������D�B��:�t���∇Fu6�(���mW7�k�y���V�k�vI��<��Bu�����tt�g�>�!2���fRp;��C-�6bl��ߒ::&�L��]����S��b��ߌ�$����L���`�%�hD33?G�M�7�	bFJBj����������.�A!í��������*����~h�����b�����������m�Њ����>��qS"��%�M'�H��_�j������(R���e0Iu!R F�C/�m��t'�1��6|��Z���|��Y< '� 䞽�R$���dţ򀢢�D����I�����a�M�=�����P���KK��|���7��(�cU;~ﱻ]`1��	�[P�	�ϊ��o5X<|�_\��2=�0GY������ ��_�?vу�D�Ff�w��R}/�������H;��&,u��S3 ��G���J:ZMͭJ؇�Ìu�#��Pn�U�mǐ	W�?��2��<5fƟx�Q�R�f�y�kU��c���-<���Yux !{��A�όÊ�/�V?�K:��d/��L�D��v �t�dN�)���Lj?�^�}eS!gY��y������Aqb�:��>��]���*��M�Xɶ��s�))��:�d:��i���d���z.�w�[�rμʈ�E��`iY��*j�{�!h�e�J��\��i�횬�X.{~^1z������b��C���`�G��\�G^}B�����6�0����{b��"O�������j$Fa�U�����k��R&d�CJH��3}�rÄO�	vl��,����~G�MQ�}�F1�-D�t�����]~B���S��X���Λ�^��R8O~�)0���َi!��Xȥ��x������Ǳ������S��J���J�o��Uz6N=�7�I/�-ކ�>��i�0���`���W(z�h�\���<�6�#�5y+��C�c���=���
4RI�ϴ�S�3G����5>Ŷ�T�9��Z
SY����%p<��M�
 �xF��]˔�!T|���h �1���q�pv��y'm��QH�W�XC r��������cl6�WjL&<�l���B:>L/J��d|�r�Zq�~��|������N~�3y6B�
��4미�(_3�Ʉg/j���]��{��<D�l�r��E�1{�7�XH�#�K�f�I�+��)�m�w72  �p�����n�%��kj2��G-$���:�a�Z��ա�9\��.nIu=�9�B|7ytrC({*5* �,0�<?�2N�����r���#���<G�9��hwtи�Ӟ�mͼ,����GH� r\�_M�9M���ckR6�W�� Q�1�@����y��`IUջ�ߛ,����^8���E�_R��1T�N*���dA�o���Z䖦���nǹm?a�K�"��w��XC��v,%x��cd��Ց{���O��;P2�����9/gN�ZE���R�j�����_��7�l<�{e^������
2�Yȁ$�O�b8�*����� e�5-��^�Ʒ ����c
�3R�Nm�)��)�@F��L�CG:��i���x�Ƽ��T�{�r�W0������Q�P��FY�޾m�#�n�L�$�(��@��$�c������;1RwO��
T�A����ӔEA���1e��C��<�C������w�F� ֶ��o%
D�$65Gy�4po~:������J5�g#��6�	�b��8��-��卙s�W���D�4���	���UZ�Cw̺�Շ���fM� ;��A=�a�����8�O7���-��cr0cT,�c#n_R�p�Y�����ᤃ٦���>3�bh�nH��7�n͊)O�!��r��Z�v,�nI_1qEj}*@Yq �X5�B��W7sWƼ:�
��zD�P�9���,�(�m�0�&��l!m���nk��|_[[JQ
2ѷ�qF]��:_�أdS��;�R�lOV(�xng�T�[�!�@\�Q�T�~��iZo�
+w�N맞�J\����&��K�O�k�fcIg1���*��Mg��[�k����mh��;�V� B~�x��'Oş�Pi^���<-�ͥl���}�I��ȿ����+�S���� q!��v�������&$]��0���Mb��a;�TY�+���b�#�(�:�q��ן��j񣭝麂G�M�I��M%A.k^P�Ɵm
y�>���ޙ.Ff�W>2��(*h$(j=�����[b��!��D�������x���� �Θ�I��� �#���{RsF�9|^���_��i\@#�
�>Q+ﱳ%��8]�p,h�(��^��&�E���Nͣ�=b���*w���n��Y��BwI�'?��S`kɳ_���~�r\_����$^�z�����K�CoA��|Y�5i��+6������~xG]j�K�8A�)�zW����@�%��]�qO�#l��b~EK���Ʃb�����~�:=AoA������r�[ �.�9�I*��,�ɚkv�hGU�v�q�	 5�4���"��V�N�B'�ۙ���rw�{}�� � ��ܕ�^ZYz���_�ɚ����z�{�uO�h�]�m���[���0��Ή��N�Q;�´�(|ӟ�bЗ��1���W�?��v߂�B�[��h�c�;<n���D��h~�R��|֣̞�K��̨ț��n>�P#����|Qo>�;cQ����.�_�0�G�݆��D�����kԬ_�����t�W��c?1!2!_m��]?f�t���� I���	#��W�өR἖.V�-�K!�(ۘ"i�솏���[�u�Db���i�:��5]B#Q�㩷�Rh�)I	����<����ˑ�����Y&�����-@��	�����S��g��Q&0��;���$�?��q.���0����G��8�F�s>��P�L��f�K"00ÁJ��뛚�o��R�����)�7�im�c>��|���K��Q�6�s�)$[u[�	��R���F���?j8o�c�dtF��*T���^N}R��c�G���zDOt��;���nh���V$�]7��Qs@:�=��=�WZkY��⭭0=�N?��o/LX�X"�"p����+�E�f��B����V�*1�_��(�cʗ��n�Q�^�) NpgY��>�wEr�)͋!��ץ�j���IѤT�왇#-� 1�y=)����3R*�P}D���s�:)�8�H�ڊB۳�/X�f3]�"��*���|uo� ���s="�G�a�xh���:-	�%�BI��}*B6C�6rU�{�<�S�È�:��*n-]=�g����K�ه۫�2�}eI��>�-E�J�ا�^��.�A����
C�o]��*7N���@��#~���o�V�(�Qk�霎?����tXlxV64EB    fa00    1f20>c�6�NYne�C/���뎧�3��'[����5n�4�t�K�@���n�r��!��)���
_K���, w;�(-CH�*W߱;=8��W>#���k�H'y�+&žO/��R,O{$�أ�Y�3A3z�VֹY�����¼|i��
�A����v�W%C��-	�'��60#][�5��˞��Zfh1���Q=��PBä]v�Q�V�P~I���EP�r�d��{=��&c�m�ṫ�3�v"���X�W��%��j^B{�D?dbԼ�&���Z��4ob��y�Iҙ�����5�f ��άn6��k�˷�������T0\$O�HC���Ь�|i/S:�T����!�QC��!���TY'�$�Ǫ��@#V�6��Z ��z����+m���/�WEo�͑�T���%jacƝ0@��T��<Y)6d^����+E'U�l�}nÓ���R=	2�g�&8��Q)�ÐDpi���2K/︝��d���=�q@�Q�>L��]o�r{��xdqw7��]uWP�g��v�S�ȭ8�\(Z�����o���O��\��Ɠ�$�9�т��Ewƶ��1a�gofKэs��xq�F����
�_�:�`�&��W�(
r�~�9\�����������N��.�/�E˪ª�m��D��Y�{q��٧#�����6�X_D�c����>o�+	�==<VF�~�d-�q�}��雎)�n����oU[�E�܍�x-^�3��8���Ĵ��kد�4��dt�0�P����Wkc"�ho�:�@/�b����XI����&n����@�W(�|�И`������k�Vg+���QAf?����&~)2�x�u�_�phh����w�3�`���hS���ˤwE��ȫ�M���c�C�]�6xOU�[�����an�>wP���t�A��qS�G}T�&H���`���Zy��y*��*�7w_��]
SvY`8ah��L��|�����7qG vE�3�䖯Hi�!���<ނz�2���d�q�z�2�0�!��Pl�L�}���՝��R�k��1s@n��ǃ��N�`�qЖRb�t�OU����5��q��u�u̅03U;߸T8�����oP�#�2�9�g��_�=���E����� ����ZH#�AZ@EI���G�n����{���:�ŗ"~u���ݫ8�/�{8n �F�`�}�F��Ό@2	1��]�=:-�KK�"e&i���~��d���g\����;눡
��\V޼�Q:2o�V?�#�P0�f�@�j����������i�k<v�
]#�>������y)V��Ay��y�d�*���8e�B�t�4BcZ����A��6t�c���rJ�xͣg��s`O��<�����8!��|p�[����e�SvX{/�RAAi|O������3�;c4��n�ٙ��^遨W�b�������2���꤅\t�����*<����Ϟ������"�{�o�;�	�|�n���?`;��B�&��F����F�{�����g��V����P{��"�|J����z��*��P�����e���;K��q��c��L`�������ˣP��;�Y� 

�G��1�E�<�ǌY�z���9�5T%�2ƶu��-��Ţ��q͗ilx9؆��'��������$�S둰�@L�N���(.�e�3���YC�#S,+�^ r�[yTJ]p���#w�*PrZ3���2t�7X?���t)�'V�$�����7?���"��m:�������G�v�%[#<�m�	�۔�a����Ǡ��=��\�;(�SF�6dRކ�֛U���E���)�
r@N��2�}l�O���J�n��w���~�p���T4�	�t�2|H.}R�H��z�^ o��Mf�R�����^�D�>o��M��lߺ�����(V��k~�ą���N���g��Ȳo�y7��E���iI�����AZ�CD������[�6Sa)���4��N��{�ɾ�Y�pՠn5�T����NO�1�C���Mi���8pd�x����qK�G''��$�2�o��׃�>�o2_��EH[����
;Z�5���f2F.Eo�5�Rͩ�T]%[�Q�R�i6*H�������Q�m��рEXǴyU���Zu�(�&6 �@4L�<
A;^����	e2�)�{k����2����8.H1�ԣ�#���L��f�&�9tuk�k�����Ll)ߕ�%y�87)�{PDQ�cG����\���A�|q͙(�_�7Ud �G��$l��#I�ܘj��,�pM3Չ�w�{�Έ.�������4�y��	"}A�<�;��0!���5�&@"���5U���G-�8�@�護�(��O��@�k�NJ�/����Vx��/a�zk���Z�G��Ng�x
���T��U�F��>�~�E�.C����h� ��	�ъmL�����a�P�aH)��Ia��jm��z�b*X��!�a�f����L���~�s.(}��!ò
N�>2��F3WZ�t��$U�6c��q�0��dQ��0ǖ�r�;�R�;8qغْD")=��v�A��E� ���~�;�ev�?ysu�	o�S�/I�&����aq>r�~9��]g�_po������v9�^B#���M�Z���9�=���)���i�3������'�4��M�S���>��
��o�����|P��*d��ކ�COa�d���cŪ�*�cx�G1�4j�m�S�-��?�Y�	�I���+�������|gJ/]϶��W�I����-�[������($u3��e��>jټ������3���g#J��E
���%n[Y��Uy�깜���m�hC|���bW��ѳ
.F�ž�89�)�έ��zl�BI^�R� G���iN�y���y��!�#b�`6����iA T)��`�om�"|�M՘�u6�7j2шY<�C7���	�n ���'�]�y �U>�E���-|��,��I*ǵ�����8�?)��_��:۵� ׎� ��7򲗜`�:���;(X��!�;�>I��A�8�U;��c��G�qC�r6��i��1A:#���	R��c�n�29�hj�����h#*,�G��̚A3�����r4ɀ�	-�Bwc��L+�%��\i�*�{@����YE��w�?�<�"e�/A
�����%�H~�-�Y�*�Ej������a��p�c#.�w�wxΆ�0$�U�H��� rtlY���.��9bbY��V��U�����*d�����>�tQokk�X-޶S=���ɂE�aNq9JY*;7(����Y��_�5,]3ܠ���捹�%^7D��K��r��J]��K���E���xlܭ&�'I�6SZ���=�[�n���Y)�o'��C)us�ض� y��td���R���h��C���N�$#��&le��W�01g�?���4�orY�f:��B�s�n������x��=�O�n�D��o�E��25$`��L	;K����_*g�*qT����Q��1:2:��
�A�5]Q��f�lT�˾h��7
�-�h��Z��G���D�MuyY�fWVI������ј�_y�W�$f H���u�=86�I6?D{�|�����> �9���v�^���X�0�LK�#��ԓ�`s4'��1�#��=��.����6P����R��椆����$�!+��}v���Y�%��JE�����`�j=���]���ܭ�X�~���`�V�I�x���w��FAGo(�\@U�YD��[8�p�b��l��̚խZ|������Ҡۄ�]K򾾂��T)�oc�Az�9��IZ���ʉ���s{���t~u_'��Ы���n�RG@��$$�.����Y;��1^��~ْ��<�|�2��̘��3ow��[Z72��;z���O�k��)��/8Ѳf�{�ie.���[&b3��@\{;�c�l�$@"3�H΋�{�&fU2�ºw~���t��� ��M n�SrV�����j��:_�:[���c���e��x;���-;�i2�'ˣF��Ơ�c��:�\�J�,Cz��k��I?j四���Av�Ò��6�IU4�[̏�`7��K?9��5���|�s{x�jڨ����,��KS֧�� P.�Iw�8+�e}������0�
̷��0l�}��n��0� �+�g�g�g��f?��zw�z�"L�v;��΅p�p|qU��Pkw^��������-�rYgg����q��Z�=��ߗ<�)cّ��~>��Xr��g	37��m�d������V9V:J��`���bb$���K�Ŋ�:U��V6T�����|L��ݻ$Wb0�������]||�2�5��ܿ��k�1�nL�&+��)�7	�c�,?������T����y3�����B�ոa��	+������Cy��+�W&�y���� �ϖe�z���!ļo���F4ƞ��C 	�al� Yfvs��C*��Q`���Z�f�tm�K6&U����?������|�`͵��!�DM�g�I��z�Ͻ���*G����ᰲ�z���WvE��W��/�B��'�--rI'n\�F2V=J��@v�9<,u~����a��P�]���#7��<͸"�VIZʢWZ��5h�7~����g����~	8���f�$�m:��'d�3��?��T��)���խ�����y%%	]��a{���������Ǣg�~'��TC"��y�ʷu=�XO�L����M��Z�������N'(,x�N�o}�l�����>H��W[A�jI��<�����ј���O�J�q�E�]���η,��-����jN9j�w��HsuA.�T��s�=����X ����Nj�l�W��@/��y�ksp<��]}��l���9�_f̗t"�.���R*�$�ӘD�TBt�_��>�I��'l��!�p�5��^8����H�=�r�X �W��g�5�A�� p&=|�؁?p(ư&�0���(6IW.Ã4��L~'w��W��Ѐ��HW$�(�lc �.N�0�U�^HU�R�(Ԑ�R'��>�� ֑�W�xA�kEhQM��0�qi"����WR���R�߂5,��u�/ZH���d�ٟ]W�MQ2�E�����v��`S��}.K 4��_�ќ��ŏ?�")#�
c�E0�H��%�e%�`��� ��JbQ se3����dYA�Ŗ3Q4����z1�o|:�,+\0�����4��uaFQ	8���X�=�^����ݮ���]́��,�L?qć��;K�s+ʣ�PHd9Im
c�fl\��H������H�IR�BR�w��E���T�����_8��'��Gw�8r�t��q��!��__�V�?I�O�qD�UJb�3K�"�RR��*��!	Q ��c�ff��J?|�ɪio��Y�
�j�	��k�DS�����- �����~�d9����xnR3��@Y=P�QC�.��\J��w���\�<P��f�W��Mc,3I7���U����$U	n�ۭ�b�����	�0�$��Ž���x,���|j����,�;�!D���@X�ߛ�V�i�5E��`����u�4��p&}�-����v�WP�<i���le]�v���*o�y����n�ƍ~������_p�By���H-h5C͙�G?	�OjT:�e��6u��I�.�e^�i�zj	R�����L)�(u��0���3D�3_���m���d|�T\�؄����(���"�O
��x��Ӭ��EO��p��
97^,9�1�ϴ�2H㻜�su \�����Q���,"��'��A��\o�+TZ��e�Z��1lhgݢ�-��&&-=��k�K��U�̐�}�BlJ�3��('ݸ� ݩJt8������5�q�[���� +':�%2�a�^l�.�},h���g�dfTrb��
�xP����E�P�a��b�����:Y��;Z(Iw�{{0��؟�gz�,�z�"c�ڟ��<5�6�@�'��3��Z�lJ�}�һ ��+<V�`)YqSͥ����{�뛉r�qX�t���%��������X���$��6C3�����ֻ�Y�c�݀s��P����Uh����Dh�i�K��/���_��Y�kݣ�q����Lmxkh�pw�1��<���A��V�o�uG{���3���]�x�hE����
�R�������ƢB�P͇�$r�+�g�E)5&�R~�P��}�������zT�\)h��'%P�1qK{w�!I��#����僥�IQ�@DOv�7��${����qzh�qDY��5�S��@��T���AY��ǡF}4A�b�%]�I�a1<��Lr�����8�xѤl�>�J�'i�͠T|��Y���Bn��Z�ߏ|a�M$e*[�g�5�jr��ԑj�]���d�<[oy�/a��;MW������-�NJ6�u6��t/� +��/��]��
�������g_�F�r��y�P��^�����aND�%�vf��Ty���ā�U��V����,"Q���[H����l�[@W�_J��4�E�5[	�Ǳ�ѝF���T��
�#�_ㄆ�
��t����o�Sp���jD�%n�,w��oy��?�Vr��ݣ�c'g�'S�.����)�Z����O����@�;G:�廁�i��Z��U�r�
��$r=~�%�5R*y@�2rU�_P9�
�D�٧��>9��Z����`��\�4ˌc�H���{����4��8*9Մ���{�4Ov#Pk?�����d2���&�J����W�	�c�򘒧���[���m���`��n8�xOC�k��O}]@��ǡ���������wH��`������	���1?eP�����Ś\O`��_��&|����&g��#�s1��O����JKo	3q>3V�	�tC{�`����~.��N����=/�؊&u1Ҽ�Ѧ��[
<@���ìP��an�cL����8��lN����=q=�B�̜7�&=��'�;����׃�v�H�!���;��ET����#��lz���f��������<*j����7xl-��`�>�V2�ŐY�:��n�@M��깆�]>�a
��;��mk�-<���L򋮀�y��[�ň��������6�N0#nD���\h����w\�e;n-��f#D�$�{#�p�>k��|���f��U��&m��r���uH4L�q�!��re�i���]n�Cm�&oሆ�Vb��E��᥌�H�����d��Qv�N�b%�&l�U!2���*�*F��	ZX�I�q��l�ؙO�0�n��7G���>�1k��6����F� ��v#+킡�h�4����2༳�����VUE�X��_�6N�� �4o+y�)M�����R���rw��C`:�7��i?eg�̰�Pe�������O����Ve�/&�������xG���>��>��OMFN��½h��+׿�R�ڢ���܈�?�J���� կ�B`��x��S�;��͟���e{Z]�nq�S�����9:=P��{���P_�_��kK���[&P�8@�B�����g�q��N�ơ��Z�a�X���WX��~Hط�>�Ev����T>oO���|%)m�C	��6���ҥ�t��P�&_mr�V'	}T��,�hI������;�M�G�����F#R������ Z�i�L�����1n��}De���O[�4���?�ɝ��J%���l����e�Iv�Y��/�#�Y����]Q���ˬG��� �����Aa�XlxV64EB    a080    11c0��-�����F�@M��-#4N��C�1�����RɈ,y=.���vd�G8}x`�&i�;�b=�Ѿ�sNj��ws>\j�_
�6��@s3'�/�Y8���b)�?��<�Q����a�:nE=~;��+$�x�b���	���JH3�������vʘ�匛"5;^��DI&������b1���;U���9U��C~
SЯo�M}��"q�k업�7�\�
3�[B��z�t1����:�ed=���	��\0}���xi
��/�#G��|�e`g��t1'�c�M�t������e^�һ��=S{f��t酔�E|���b[5��{U��\���c^�̅͏���tQ=x�OP.r��/�CM!�w��κ[/�}�>��pI�w�r.�SYW��W���?�ꥋz-����YZ�����x��-Ͱ�Zi+
�����Y/�������W�+jĘ�czJ����<!�����g|3Uܻ?n�$��	��. r�P4
Դ,
XGYb95�>�	���$���g�s�С�B�v��cсI�y1���i`I:n0u��g�\R���ցy�ĥL�����D�ˡ�u�uj��4�<2�U�T�U$�J�uY�1��ߴa��VI��JE���R��J���q��e\���ٺb7�e������������
N_'�f'��Ch�e�U��l��S�T��eh���>_�R�N��ʊ�5B?¤���M4�����J�H�,������plJ"ң��9�ʑ�E�OtQ�_~�d|��a�͖�$��W�6N|���1�N��*jٍ��Plȉ�<,X����?w#�vc�����1�s�����m� �}������"�?�s�rݶi�cx��ڃ�5bd����Ӽ�B}��1cRM���f���Y*�� G�ZX)�?~凲�N�Ar���a0��b��J�7f&���*+�����RY�\�vaT�u
bYZ ����b�4Hv�e�!�gm�P�������<�� s֥��3$��r�NB�;��n��	"Y���N�HE��lrMw(�ٜ.6�~n�� �RlG�tLU���X�����cڰ��I���<�҄��ԫ ���^>�����#�C����-�\��'$L�X�i���a�q�.���Ebp��+��*@x#��O)��A#�]�ZK��%e]����BC)J�ы�6ט��J���C����d����5 ��88>���֪�6�kS�*#�^��\�Y��䔎r���e�)��G�p�)���2�W�����n��[��@Q1VB�=]����8E a��N� �Z��,92���=�P�7��m'Қ�귙x��k?Y�u�F�y������ �_+�z��;�6�o��M�(J��R������E۰cd�ѕV��i��*�o:��b��p^s���7&�jS����#�l=���%�Io�<��)">�,��v?��9�3'�ȭ0nZ��g��k��E
̐7G��NJ?x���+5u:Ρ��r�~�pJ",œ��&닣h8�pe(�G>�;��d�N�?�r��R�ڄ�gv1 ���vsT���2��j������5W]Η��%
��̵ET���b�:�'c��p�[�.Ԡ���x���!����X\�m(��H��׈e-]�+�q "�5�
�sҨZ�S�e�_�!��±��/.�>���׳��n����.v������vK'D�'L	�Y���F[J8��W��2ѭ� e�'��Y��!�#�gP`�t^�g\v֕�f�z�.��[���au{J�`�ۘ+.��<�ӋWE	?������/%ǂ7��u<AX�ɦ!z��o9�|�;^h��?���B#) Xo4�W�qM"�Q�P��+�J�6�������k��ZZ�ܔ��.����b��P�LҫH[�2��Q���,뼜b���S�p��h���=�0ئ�R��~o��� ��FK`ȳ@Bսz��m	��Z��<�Ɠ�[�0���l�]�H������W�
sZa�IAF�K	��I�ҵ������]/5ɤ5�,��,
��6���i��*N5�GCE��k�~%0��u�rA:�����
ʿ"(��#����B��r�Pb��(ؖңg�Кw�:�� �cS2�y�����j��/$~c��Fm�O���=�k2F��j0!�5��n���\��/�����K���U!W�y�w���MeH�9B�t���s�%��/&Lgp���@���l��$a�v��r���HܢG��r�@u�UgŌ��1\K�8�Ws8�����1i�uI62�y�h��d��6�Aܹ ~uK�z���ߵ�ZtB�vi.�� �|�VQ=Ɛē��I��%Yo��2@ ��݊Q`�J	�2�|�1����a���p}Y�Y���j2����1&��!5���ce��'"=�q_j��~�γ�f�
ȯ���=�rD���RXF�^��w����,���U|[D���y��e��)� ~B�<p�At(�f{[�ȯ
�[�hQ�Tx��mM�bR��Ě�:z'xg0��cBc������;5/��}�����J~��~���Z飩��6�����b�*g`%%<�n��-w8�t��_ߕ!w�L�0�`�-�a�g�m�_�Y�TX^¤��7�tIb9�)4��
�r8t��M׃��w�K�f��V��I����=�-�ߙ:�G��Y�w��/�}�%ɘ,�3�ԇ�X�FwY"�ȡ1��FcZ�t�k��|'&w�Mct��痬��'ƽ�T��s�|l@1GI�JV��l6��`^Q{��r�kNH�RB�>�ÿ��\��lQȽJ���M\�k1�l�9��ڄ�Z�Ш�Χ����۟�����z��㫙��E���&��Ӗi�>�+=}�'W>��W�B��z�Y���Q�o#QϘu�knxO)£�媮�><�F�=_E�s'��>i^d&/� �MV�Y8k�}���L�x�� �@x{��j� �_�^�S�d\m7��j�v�av���:B9'�ɵ�;S�.gTX�Mcq�	�P�I��U$� o���[;�Ե>擽#�������^72�:k�Ow׸�3�d;!F, _(g����T��S�Gj�/*���?-Oب�q̹�',����=�?ǻ���C6z�C)٭:^h< �q�]�[�Lz�O�1\�D?>NHa5S�
V$�.gkW�ao7��n����oR�cU8{�)9�v���}0K}XQ�T��c���λ6��#�8M�$?�/�^9���^a�Ud�� ��� y�����Gr��@Z�bs0���Hd����YDjvk���mb-I�?6�1>��װ�U����%�j�t����,NP!��l�^"��8�����_�~ݙ$�c����؄�ьB8��|ܸ���G�GG�R��Ȏ����jT-x�?�q2B���9#=�=��ݺ�4��i调��[���|b��XF������=d��H�Q~�8M�\� lT;���fb�#ŐG�8El['H�&������?6qH�.�ק���%l��K�8��ܕS8ֆ8.po��PH�.�%��qʼ|���ju\��d�i�Z9]��E��ᨱ:E�4c��h��V]�RE����'�}���x0T��ف#_�wh�޹��+��/*?��DF9�#a��p�P,��tӂ����g�[���9��W.|�ݤ��X`@��6#CA���B��*� ��b��xh��7'�MU>��gG�|����Xr�v@���ӛi�B�f�8>lD��;f�B��6G�]�#ޓm:�X���yِ��
-:�Ӷ��x]��I�ɯ�	:�0J�PYpnq=����b���V QhU�P4:kn\��XU��z:�Z�R�x�G��HͶ������=�S �x��`�A�L���%#�Q�p@=*����e=p�!��jz&<]B;���[�(���]uí�)���Bbߓ����\���f�]�  ū����G� ��8�z�Ñ,Z#K���7��
|��*��i���wr�o�!�.'�1�2���V���?���m��[4eoD��'VX��l�Z���!"��fK�"��$�/���9�2b�'���V�������)�f��Z�^H1� a+�{�!q���H��ۈrt��'R��QX�0g�k3LL�Ʋ�j�اcKJu T49��)r�s2����N�Tik.|㉻-dFU'�J��QⓌ�!yƂ3_.�q��f��|=�c��[Mm[���p
�r�:Įᔶ�[s�����������Ed4���Qd���FR<�u�c%��U��=�f�4��S!�i���e�:�ְBDGl	2�ϯm^�>O�}$���g�a�c�Au�l�ES�A"A=-��y��,�\��c9|���Y��hRv#����� cs�OhG���X�릛�ֿn�����0#�URV���6���uCG]s