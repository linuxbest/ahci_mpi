XlxV64EB    fa00    2e20�d;�<��Y3j�r0�x��/�P��p~0��Z�d�eH��LiPJ�)����qM�;�]D�)���{���7}���O@"�����0ȅ`���EX�0G�T�{�K�v������'%�0��g�|���VuJ�[�hͮs�B,��I� a��/�L��������G��x�z�����M�Q�戞�2?I��l ��_O�A#��4�6d��
I�b���=�5�aq�h}z�����)�z��(&�	��m�����A��!8߲Q�_-o~)�1M�G�3��ӶIZ$Dvk�d�K� ��&a�:v*�S�)�t,3���؛�}<�O����K��e��X����e��?K9�D[���G��ӦK���U�Q��m��S�<�3�a��mǇW�U����+�"،j7����u*Z~�,��gC�����?7�UJ�@ I/�_��/�_v�������sG	՚:���8R��1V��ߥY�������?�*����2l�*��Gl���j�j��
ȫi�:�"�P6w��~�7���V:����s9h���@��.pc' HDT|
�����jK$���rڷ�/i��%�?��V�:�K�W.���8-չ;�o�~�h9IV�,c{O��ݥ���A79�MZ�J���4Mv��˸���+X'QWa/�RPO.�>�S�c��m"�
1�FN��U���^�l��F�4h.`f��#_+�2�ًf�=#ܬ�P���d	f��"Y�P�ٮ��F��o�s9u���	���U+�c�b{������li���`��s1����=����pb8i���,�hvw�t/"��,+� �'`Ň�i7�����p��p�����!Wh/T�4���S�W�-tb�Cr?oK�*
vY�l�wD�/
H����w$84�����;Ed<+4h�e�)�N����}���p�v�|�6i�E�ذ�+'Gz�S�Ԥ~�oΚo��c�.��(�W� �� y�VƟ���K%<{�VÆ�t��r��u����	�̍� 3�,��u�4���se����gB;���*��+R@7p���Js񞛜p�g�a�{��ց�D�XyX����$O-gn#h:���X;�����.Lx���'�������Z#3e3U���̰�=�T}C/Ƭ��#̪5H	:�mt
 �	~�Dbҗq�$#$�R<	Sȥ�@B��=
��c
0mA��Ǘ�k1�,&k���~Qpv5}qL�ABurP���ao�̿�����q�|ᨅyh���U�B�|�!�U!�݃����!.S[�����}n��a.~τ;.uv�q�Mr�����dx3��AungbS�X� ��&�<���o<�솗j����ԇ���ɇ�S��rb핹�XX�o��7��H)����x���T��Q��A���X^ϸn=jS=m��d���x�3���(h�$���찝?O�cT�P�^��S>����
]k� �g�t=UNG�
����f�>��V��s�" ���������I`0���d��`��5�X�V>q2?e8��g�h�Y� K��$ؖ���m�O(`y��q��~X|�ѹ���� dS��AP_ZVma(]���b]C���})^H�Qjm���#]�ӇE1&-~ו�9�����䣶��/�a�b�L�d��٦���D���R
���� ���"kr�4M��Q�N��	�b��n�(�2�3�?_�{�p������"6�����Ikو��Z��ᚊ����Ee҆�%�yeU���S�kNU��6�$���7�qG���[o�ો�N�g����j�@���-�S4�r)3N�$R�2RܿC�"(�Ar��貈�����ҟ�u	b���M�6����]������quW�\���<ry��#9�^ ���+�j�ٜ�;�@�MZ�ط�耭B��z��mA��ի
�H�du��8����弜-j|Ԧ�'���R������6#ky��	���uM�����~��5	 ���0 �S(:k��
=��OA硵~7lp@�1�צ7W����-$g)Xd��H^���:*ô�
A�9e�.M��7Fm�˰�v�g�ɏ��I�2!o����m��q�{
ܡ��k�b]O���Y�6���T�ySG�D��5L-�*J5��ݎA˒�~N�Pq��-V!�Z���k6�	����}��w��_�����wQ�U?��m&Ev�u��(�=��J*���7����z�A�4r��*�qI�!kK��Y{'֖� ��}6�{ŕͅE��ow�Syr�)'�u���_{���j1]*r�T/
�;�&_�K�/y�LQ޻�B�"B�vz�C.y8Q�ǦX"�O�hM� �7�"��@�������v㈼2d0�P��i#����,��rv褗9w`z���̦y���Ё�w|��tn÷�~���8��ÎPl�Ә��Іʻ�G)~��?���s�W������!q��0^��-�]�Io��a�ݼ͟��gÌ�?�	3�c��r�j�>�F��ߠf��1t�n�
\rf(�X��!e�8�C��������ЃZ^��A<���_6p�ð��1�X��� r|`hB�<��k�\���kI��sK+�	dt��	bb>�`u�f�7n[�9�C䛇�&��\���H�6�����ɸ��\��?3�8Y�F$y̽�u�5g�%�Ѝ%8�D\��y	�o�ڡ���z� �n����n�xU�dJl�"�C���>����,�86��n����:\e�r��M
�P��=$\���j�M��2�jY�_��ߦ�?#����R����Nۉ����o�@D��"�9����
��3��n1c������I$z��¢���.$�E�4lU�w�/�ׄ~��7�[�'?o�>��nxE�t����a@̺F5o�n��v�B���+<ύ���19	���hy~SƱY�|��%�{7���J���c��=ϛ�cm���XY��� E�r�="�	DN����fa�X����@��=��Gu��s wim�]eu_̭5d(j���F��%Z���?T�5�_��I�'�x�`,͚Π�@���].������"B��ԇ���Y�yP�ke�*+*k�H��nI��1���pV=���i��[-��*_KQ��|��(R�^��r1e�*@��
=F�� ˎ*�P�hs[u�}�*�Oo2�I{q�Թ\�#�Fứ!��-P�x�3�uK]��+-U�OsuԵr'	׎���?�/2���CE�.����ckn����LP��<GsY~��3ᓮ���*���]��ɵQ�D+a�NڵR	*�40>����z�+SӺaI���5��"�T�"����:k���z��i���Ns�R�!��|TV���V1x�5�h9O�wb&�����Յ��Y�������z]0�W��H�O8g��	bb�ecfW4�F��i��)A*��nd�W yf�M�l��Zҵl�yc��q�⯥���BN��R؀�7*P��@u��`�1%-p�y}��Yb���B�`����1���V�81;�#xb�׀�yy�Q�wsǐ^��{R�� �~���F�!�MZ^�q�A�mۖH�o�Uo+�x��ӓ��K@���E9���c6ל��ݔ��ƹ(>�M\�I�]�9���P�,IFqg�t��O�$�)�l#�ت驞�BE
a�A^�~��.�fb���p�X��%��`�/D�?M8w^�NU�?Zխ<�,T��U'��#�w��rέ�.ҕ��I�����֞�K�+�nd��J����=����9>�\ˉG�g��q���j8Y%[��}M q�h��6�I���]�ڭ� ��� }!�_!Ht�|�7���_D�Ѥ�Ji�ь)9ǇN.�3sGY��Ț��/td�\����zڂ �ƿ~B9=�zH�$�kj5?�IMp] ��Z�r��u�6|d���=�(���%�#+��s���j56�Cr��2�\��)	�t,��CS �$��K(�!$����q���1�E�%x��F�Oo{F���؟������?t���D�p�����92���yA�c4[c��C~�o�q_�֞���ڨ����Q����ON�҈}�����pZ�0#��)\��U�2�ɳ��!EQ�XO�$>Y����S;_�J����uz��#���E�������M��K�i-P��m���d��S�XE� N~��r����R�e���-1Ѭ���M�3�.���
9���](-�������Z��!O!vZ��� t����Q!�de���oSi�IQ�tr2g�'A�=R\Af�Qc/�+A]O싪^��"{M����M���cb�	�92< c��-��م�� 
�"��a)$�W��Ȇ��!�V-I+e ��.ڝ���c�~^�C���p^�R��]��č��J��� pnk�=-JA��n4��<��}-��2�QbRţ:��L�,���i,��Yq��u�f�8녅��Ŵ������d�Eѐx�=��.-i�;��m_\f��F�q!u8I5c�~�/N[{Gi�y� ,� �������|�-5�#����ӹ�F��4��Y�6Y맛�IJ?Ƣ�����t	��)D����cB�L8�pي�x2�����b��o3`q���l���¾��v�£��z��'g	S��ZXC�V���Vt�Ό2y����p��b�c|�K����C��`�7�cb���ާ�,վ�c��[����D����C����4"&>�fj���t�;�t��*U�=U�wo��P`Ʈ����C!y���>�W�XϜTM�Iy<f���y�,�Q��$.�Eli�%��/e��� ˽��ʋ�G���>�a��qF�Ʌ�SY�rg�IM���#�w2cj�t�IY^��[&��:2�!���%��	��"���U�r�����>����;Π��0Y��/m�7��z�AW1je�a4�n��
n�ʜ���ݫr���\K̼�t8����_�#�|D�8�f�\n
� qݞ��3��"��K4IkV��u�n�4 ���>_|�� ���i�	�a(��䰇''�G6S�o�)}�!�=L�}~�p�d
~uF�/%F�e�vE��fH4� 8z	�ݞj׹ms��Hz�cU�J�o�ő;�~�j��X�:N�򋭪Z�$*-�2h���/[�'
�>��ٷ��Jč`�-�1��z�$���r'S?-�:����B}d$靥WPP�����fU�s
2�F�<��<��v|k�]�ρ�)fwK�W8~Ɛ�#�T4��'���_��lk�3G���S��Ѫ��V��9��TJ6΋��|cڡ������㲟������5����O=�Z����a75\����� �0#��WKV�wƨ�z����%,�n�,�n�m��$��θ��3�����LWO��KXC���$y�C��]z�^:Dm,C�#;�B}2~�y*ˡ�:	6ޞ �w%�x)g����H����\g3Kvֲ��xeM���QC؏,���@�M �����ʜ��w�0;��u���2K��ҡ��0��G���c	�.�uqd�U�`u�Lv.i�����r��V[Y�$��B3���[��X�n߶�7��I������{�+��"ۑ?���8[d/^�Nk��u��	���DZ���@�O7��W����n����ϐ�A1��gθ����q��wx������r.��
_�r�c^g�"�r�vb��l�m�=�����=9�z��ښP�9vD�m�g�����[��R`���B}�l��S�7!�~�/�Ӥu�ɋ
�?�.Ap���Y��)�@�YX}^�����#���W�4�S��P�����?n���M����8N謗���TysY�q7^ю.���T�Y�A���=��&v�픾ߎ���=�{�Z�^��E�ƝZ�ډW�P�=��P�bm��W͆.�D��v�7��Y$SE���l�5�]�όRjf���{O��� t��m0ra����v��݋'���x�֮�ɥ �m��d{�ܨ7������]�4�D�����Y_�1���s��q���_ȳ�Db�����<�z�JB�و�#WVIfe'u���mfN���nŘG�B38%����炰Rr\ą&����5&ߥ�;��.Τ�w��_CY(�~�G��<XPbm�8�&�f��qT[x�+��*x�Q���-��$��Xz��ۉ1���Z��`��i��:��=�ªјU:6��M坨h� cP��:z6{�}+< �W@�� f���t>��+4���JL����2�ѩ��I���U��&z�^�NA�5Ҳc]@�UY;�U|�$+8�{*_���CN;�@��o�b���ɬ��9��5�_Xs�d�����|�!�yd�A�,�Ӄ����Q�[����]�x����J.�C�|�:�Ҵ�2 �Xa��k��V!���|c��݊VޏQH��vv�5�� 3fIGV^����#7B:J��� r������	POM�̸w�j yl���&�����9�6���λ�A
Y�*���ُ�����{�l,4n���)z��Dn���/$p�A|�H��-�d;BE���B�F]<�J�d��"��@]��`��LlV���gkH=n�J#���$�����K���i��#e�n?!�n`ѫ�t,�턕���^MA�J���h�9uIgq��l��5�/�ޜ3���vKRg�h�!��(���"�ma�&��'H���}��Y�v�]*��sV�żt�H6�~;V�����R�� ��_`g��Io�s�.UO�5��0o�YY�N����ՙ��6��
%���B�P⭱g�W�adކJ��\���Y�[�P��;�"�C��Ԛ��S.uzd9�Ѣ���ܖ=V���w���$�dD�d,9��h+M٠~�|�"b�\�!ZVRP�>7��V�|w:�XQ�����4Q�cC���B�^�nS�z��i�v��1JH�<�(��U������e��?E��,�v�Y/����ߠ�Z*P
շ��Z�s�qm!��;�������Bop�����M]:Y�w�����S�-l���{��p	dTc�y���Nbv*��pec?k#ܸ�T9�ٮ�(7@bX��|�Jz�ՍN�X��Pрe�%��W*��׮��=�I�E,�Kfx�sҝˀ��~F��uTp�
V,�� �T�*�mlc>���ߢ�ʅ������m�D����l��م�s���3��C'1+%;�6��?�?�Q��v��b%�/���04m�Dk�_ڍ��#2JOB�����d�����H����E*ͶR�PC3O?�$���qy�����Z��`���a���4����w��B���ǫ�(���w]�A���Q�i(����\�"ȸ�u�"�X+�/?D�)�Κcx6`��r�L�i���!�)b���"�Z�(���u�m�a�.��eq̂���R.i�@�)Bh⪃ �z�����lV{��+����ݙb���y�k$���a�P� �/°��󊋗��ڛ�.�͙A�>�PI/.h�SD�_�|�����:,���U�	Dk$�]�;t)�e\YS�
yf�V�������]1�p�P�>��a�-F��*��Ks!i0s�A~`N؃���'ƶaYin�%�p�N�RN�h7q���P��HW��ݟ��l��Sa+l�x�^+�y*w������ma�VZC8�/����z�.�s���Tq��` ��/�V�~���k�%��Cޙ�*�Ba���	���'��85���CڲF�����$|�� W��!0�1���5l3z�{���K�|�Y�7O w���]���-�UK��p��g}rΨ�ep�D�`I`�y�w���B�i"u��z±������F����P�ԵM�LU���������ۆ�al���ӆ_C���+ mڐ�����jk���WIѹ��a._�;t@6�����Ш\�"��m�^;�t����YvB��}�u3�W�:
���݅�����!}�~���gJ�o�b%"l���)�/�ۛ��[�sREܥA�Xz|�:a�$��z}�hx<����4L(�[.���<��WK�jcnB�``�!�����{��m^�Vo�Up!;�����C�_7<�=5����~�����p��79׃B(���b�uR8������qS���Y֏�[��u�+n��!\W��.*���XW��m0��-�	�=�,W��$�#ۂ4���6���B�]F�8�J�w?��*��0����J�ؾ��2��E�y��MQg�*=������2�q�\
Po^{?��.�#�(]��8Ipٵ$�ٿ{Y8|�>]�������S�!�ꎪ���CY �#���dK+9Rb:&#i���9f�9Ni7z��*�|itxdH5 [Y�+̞%������]��=�� ���V�l*.9@�"�DD�����O�+݅� WMAh�7ma6 x�Xu�$#^�s�Lã�*�X�U�D(T��:��Q��
���C��Y��`Ms�-塍��6U�~Z��֐2
�HU���F*��[<���;��V���7H�*C	@;��G�h&Eǻ]��dG؋=��NS���P5n�H\N�̵�1�+���qv۠M+h��v�^Ǌ���zj���)��Sw� ͆��5r@d�MLyD�c��]��S�2OsRv�/1,�vš'�+��0}z�4֌���,�|��.��W�W(��k�|��/vm���0�G���.�������f2Y�v�G�	Nף�_ӏ���������:wt�bw�ґ."�C��Y�����,��(��w����>ӫe��%L>�K�E��,2�����nui�lZ��y��z�l�+b?�_ޓo�{��l�%���:3r��~-��{)&M	��1���>Oy�7��2�����^3_�$V�yOd��K"���	,ͭĉ��}nN���e+ٳ�����ݸ1�Cظ �����b�[O�����<kYC+���C�>}%<�1���61�1Nj[@��i�K�S����S�\�o��]�<�p��:��<ǈL�[���L�-�M�T��u?� ]�r�j��F��Q�%8v5nզx�)�@O��$�}i7�,:S�ᯃ�U3�5K�}�����W�vК��8����4N'��uJ:@�e��U=�4(:�>f����`yD7���>���!�/�������l��ԇ�Ҹ�s�QӚk��󇏔��;p���Hb�j����s)�h�E�D�4li}6�d�����Yo}k.M��}o�D[�U33d�(�!wl��kx3GW��Ӣ�+4��	3�L���,�"��󏨨�b�(�>���c�4{:�NB �iפ�	.9D��6�9��!�!}2�g��̓���c�$8�St��Q�Va�B1Đn���X�o�(w>�ץ	�kU�.8�r=�Ha��.R5�Y�Y����ҋ�M�lJy����c��[>��*61G����t�+lԃ�6j�+��a�#ϑ�Y٣��a_~b��3�s�~ �镮�����wd�{�*W�� ��٠m�YˈiW�T�[�5�M}ލ�T�>sH��%������%\`�@0��vq�d�.�j����s��3q��.>~��%�<:�I�����ݽ��e�n����]uw�0�*��n�
�},_�&���2�!;�E�����'�+hȾ�gM�zɮp��_`AfI}.�����7�a��Y�l�B�SwRc�M�I3a�i���4����rh��0$I�����u��P���B�ˎ�WBX�X�Z߻�,f^�vZ��}p�b�n=:�᧲N�-�j$�-�!���E��.�����ePa mҋ|W�>I9Ѝ��G���kS�{���� �L�>����c�ل��[� ����d/t1�)"	���4-��9���o5s(��P�r��k���`���Vi4wӠ���+���F��~ԅ`�l�m� t��&pm0�%F/P�av��%�ɬQ}3��	�^M��)e3&�|�E��c��.��/ѬG��mFs3n@��u�<��SH���o���Fs#�qW�cFh�K�&k�=l���f�o�9�>o�EF�Oi+0�Qԅr���%yIT��ɔm�0�OqH�/5��6��5=ea�$Z̠��ś�q����v�;��,�_#�w[�w׾i���{�t���k�5� JD�ʋb+!��y� �ݤ�|���e��k�?6Á�)yl����Ut��Z�����1��Uj1CS�D�/Ez$�1�G<�[���a�|�(z(�`y_���@`�b�k�B�Z4�>y-m�+�U��N"X�<��5��^�²!<y�S�w4�h�y#4��Z*��@xe��k�'�M�@!2H��LE��$ Oa���?XI@F�t�j�V�C)��a�~K����C�
���kaL�~&#�ʂ;�QW�����n��3n��$��)RI�y�1Ne�\!w�_�����a��R%�+� D�Ʉ��ܐ=K!��S_�tj�B/�m�W�&�+��z@�۫YQ�Xo�ѧ��E����2�#��_W���ZxM�H&'s�u&�cL�4!6�9�ġ�A��gʽsm�lw��)�j;g��%<��!��G�tA��:n����&6x���zZ��v H肙��d�p7y����M�p(�k�����7�j�
4O(Xq� ���(�rir�TC��F���O�ݑ| ��R����6������R�}/KI ��S�û)9�U�b�U=]�8MWz):G[x0L�!q��Yv7�W���		���
30��L�yW�n&{+�.[������m���Z:�(�J��}	'�Økh�����=���_J꧇�t0v��G4���	��q�f��>�4��+�����y��!�H�� ���^���|3�=�K����f��=;N*P�;������%�����U�=�'�T��E-���}Dܿ/R;Y)��q��hv�P��F�'�j�Q�!��}g������'��@Tj~$�P�Q|X��zAc@��l"A7��G���6`����bޓu�Q.$�2�4Yb\������],��)�)�Y�%�[�����^�_�����w�_����٪��'�3�2zëe �2�Y	��������O�]b���r�O����U��'E��Y�O����#��Q�<H�2��ŉT�}v�[�}�a���ߌ��ʟ�zz J?�]��	�����<��+x�\i���*�V�Y�H@�2���2��N����G�Y_A�6����"�
��B<E��U��|�������^{>����G�3��봸��$�ѓ�����Ȧ60�f�����'nNE�W	��+��4���'���@�\��l2�RZp=�|�e|
nF�"0�6pm�q��Lߒ�,Ī6?�j6��Q҃i�5��,P�=aR�wۆ��+�RO[K��|?BJ(O��D�P+]3�,�*��,�b�JB��ȡ:u᪙��m
�5O�3E�h���I�d3�eR�GaZm����̣q�Dg��d����u�4�꘡��g����[�Rc��X�d# �q>Nb�����C�Ɵ��R˴n���k�A����� ��j�l�XlxV64EB    b56c    1ba0�Tsm������cv.*j��b�����Å[�|���5[ek��/ H�4��M7�'��l�?g�1�����1Sk�]4@���������e��wyv�;X.1B���E�S�
E��0#���M=O�ۡ��	���buX�r�?m:@��U��D�+�gρwf���M?�7g���!���=_�@���'��q�97�I�AߔfT,?C�Z�V��8�cہW���Nb���툡�8f�<���%r��1�hɨ�,���In�'�\�$V�O0#�-;��(pm�>m�k���z�,�a�� ˽
���avL3�jـ� ֈ�y��%�C�td0�	]NMިk�b��5Vy���Ӱ�=�3��;ye�b��"K'/����J���~ Ւ�q�1�M�]^���/�%߅|xa;��O��%���XL��ƣ��J�<ú�7�c�We�?�6@�^�E���W[w^�|dR��,�e��p�ߜ3�����7�9���z�M��.je&��FތV��SD�u�u\ TV���>դ9r�욢}J�����b=����>�|�1\�$�T�V�����oL�yE���Dc���0���U�e�QC�&W3��?֕�K����%s.%��0�[������PޯX!��,ߪ[d�D`_��A��G�A)�A���[()��Ŧ��L>Uȗ�̌v����D��&�wxYC��"�D��Z ��o��8�4�]3�Y3>���Ms�f�2���m%�8�{��^9��Ѥ2�V?����e��ŧw��X�"��&.j��rJK�5����6�<?pz	�0��N�|�et$�u��Z����Ɯ�f�4\�G`�B�cNv-@y�� $x�VZ�i���m���eO�J�����nB���0�K�e��5mJ2�6i��RF���E*+�%k�i���-���(�_H<�c��7��w8P��ϷS�(+�z�ܜ�X�t�I�*M����=}#�я_("��_2�`��EY+o3v׼Wb�F�(%��34�P�w��>k��ٰoOb�,�*��E�0�`%��L�
.�?�:j,&�zC���������i�PAA��z�LL�Δ_m�Tn�%>�y���*�߇<���X4 �x,#�T*pD��������rsִ)�}�p�B�cwҼ̢�գ�RV�Nj�(�V0��h���7i؞��Q �VG�!aG�=�^�:5*��hq2�k���c qL���I��y:���	^�"Q���Ƽ���d��Q;����o?�!�,w	��(�̷�/�F�kc�vJz\uB?���%|,�3�g��%d�$>��z����A����Z*T)<���
��Wi��~��XO�Xu9���R���Th~���%�H};;Y6�����V��W�n5=��|�$g=�f�b��8:�F�����l�v �t��+�ieFo����׉%���O�LV�a"���  U�/S\�\3��˱xlGol����]���w��z�$�kc�}�&�H��jxwpMS�'ɬūi��T/s����7����i�P��N�j�F7������`i�C�Җ}���5��d� ����J�ѥUW�2aW��9-�K���c��y��)�����F:�1��GAַ��m��rp��O�\٬5I�@
q�{:�(�5��~�;gTI��ƍh�kG�.�La̐����-�\1��N��)��C�b�!�E�q�A~%-���v�Ņ�]��v����`X�y�2�N�R�F��@�8�X�O"�ڹE(�8�����C�(�Ë�]A�;�ߖϫ��,��A^���"׽[e���?#����ںNs�`�ؚ�qT������ܻ�/����پa�0Ia�cǽ�0�|��;, ;y��ԩ�N=\r\�dv.a,��E�p1�FdQDS�­�%��o��
���V���5RM ��A,N3�w=�1�MԘ��\s��b�$UD���=�'@���i�.|���ɿ]DG��z���+��R��|�U�J��Y���Ì6|�u����O�b��d.�@�sY5f�����|��o��S����a�-�}���@m,�1��1�̣��-GX ���0
�O�r��PobX�'���u�6�'���I���]`�P�ۋ:�E���/Z�w<e��M�=�\5��.�"�6T��}�U�@s�F�Zto,ȅ��A��
,">ixC��_[��.��Y�"�ɠ���є�[�������/L�����9Nu��c�$��r�Y��FȎ_�E~�q�bH�/��Փ%�����')�N%탒s�j��K��k��l�۬0�y�������2�X��s~E�;[B���zy��N�"r2��	����7�R�����(��չ(\F��x�=4&�t�|x\�s[�jG�K�R��\fU������dy���Ԭ�=��� �Д��9t��E�)Oc�[�k/�n�W�����wf�P�v;A�Io��M���z>S�����!��T�����	f�R�k�'�ݷc'�� {�73�\E�e���L�ZS������#�u܆a�@j70�^�ȝfb(��L� ��
R? 㜟sݡ�����.薐�ᓡ�����ȳ�3Vd2���
��Al��Iڐ��~�T�4nֳ2�j��K�9��;T8r����l4�0T.�FD�i�o'����ʈf��Z~#x�*gv���y�5O*��eߊ�k�xB�A �~R�'xf�~P�2�s�����G�5Fg*<XLF�5�8f�w�K����P;+�5��EO�ç#�Pk/��r��.��.23��hlP�j�2
�m��\ٟ��AF����c��='��	׉����R+�^�d�l�D��"��%��*��iʘ�I�x��D���� ��!�������7l�H�����y[�U��Z�Uʑ��ǊMS/�t�?��,�6���%�񑓩+�r����&������B��(a���$��C�Ig��G,����!o���,���up��X�� �tNc�:�o#��Fd��IT�~�S�=4HI���|��5&;�#��*�"'��`.��B�n�}b�4mXP�<����YR4.��r-��}�n|"����&v�%2�,�[�ˑ����\a�i]ԝZ���uVC�y�'h�D���[zF
h��
`��4H���&/��f���J��V���9�'�? �wƀ�"��oi9�Z�"q�-9�x��h~B>A���@[���+��n� ��N���6 Kq>���"Ã�W���Kk���'��\�(V�}�A	�Z��c~�ڔ�2����/Ds� e�w�1��Ԫ�e`P�&e���@j�;_;¼E��=?UFƢir<4	J�ǯ�A��
v�]�^�+㵭�y��A��}x�|�Ƀ�x~��SF5i�	���|��+FN�?b&��m�lDu�Rq�DzÊ}Ѯ:���~]��N��F�i��k���}ߍ;�/�_e䐁��#�4[�K�AH��U�aԷ:���=�=��K����g��ȦsW1܆���gT���܅�T��J��*$y����!���cF	��^y�Y�ϗt'N�y�/o�<�zl�޼�ݮdE���8[��[����W� �;:SX
��<ƙ��&gŠ���U�#�XJ[��h��t�g_�i�R-�Ur7�9On���=�& �Yz�0':U��i7�v����y���"�k1��=�n��O����At#@�?��֩_�Z�_��N��$���^�tWY���-�$Z@i�9�	;7�?� *��9<����X��s��k�kv�c��	�2Ma����M�0z�mV7�� � ^w�l�?��Y����JO�}ҁ����L�%m����H�#Zhqu�C{���N�{��:�d�����	�8fl'�l�{�G"!�NL�\��~���#J�)�C�[������0˿����{B�����Ps������Ⱦ���\4�1X�#ب=�\�rh���?�*d`�!�:Hv�/6�#�;O({�T��w��/��6q���AE�Q<��� ��"A�^��8���¡�x�G��l��7��^#���F3���<�����'������W_`S��l���)mŁ�у�6���;a�*05@D�LJh��AF�f�x>��@cޱF~��CW��@��/e���%������7<�J8�S�Ц��bFƱ��� ���u=��{������_���B�R�"�)���nB��d�}W�p#{�c��7��kG�;�ks�G ��;�ň���mY\a�fL�B�J�����֍*�����?����i6Hy�Z������i�u7n�X"ced��B-b�G$�nJ4��z�d���h�Fn�ȵu>?4��V�n{��S�hړŃ�p�YJs���g�;�~p�:n]Xv�S#����G��e�6�+Y��_>7L�x�mP;T�ɄA�>�h{ʹ��)i�D-��ön�д�E��M�����۸REZ_#r��#-��ފ����v(m��J��(�A9�4��xt�˧J��S�5iy� 0S��O0Xi^�8P���9�M6�{]N�Y�&��i|*2�[i;���|�*�4���wY�pIc%t\�>�}��f����cqĂb�ɇ�d��X���şhP�7�x���D�r`Q��5������+�w�����m謼W+%�����5lO�
���)w�HN9j1���b��_�E(~�y2,��#�EZ�_|q>�G��LB�5��6�ݼ(n�m����@:�8eI{��Ft��4�YUZMTe�zP<��i��nr-�쎵���y�pĝ������Q3-G#� ��Wr�+��l�;��7�hv��!�����C5c;�Q6:�������M��A$ڈ�*Db�lG�������㌗zC6�RD�Ou�8Wi��8]����7tfk1�"�����r_N����8,f���P/���B����k� ��B'���}�Q6��e�݋����oBޞ�-x]O�+T�(~O���q�T�B��zr/�Ŏ����Rt��#�Q��]���r�͠��������n�-��b3g����րl�z�ZC��K�3��'�ˉZ��D{&������WX�oQ�W��G�tC"�IH
�eT ����/�,�X�lW����X`h�Q�����z�F� D*���*���`����N�^���qH `GvCa�?^N`�"̧�.����3B.NL�/�=Q��o�N�������&Tm;�L�8)�B�K�p�ps��HS�jM�9d0�FyN��^�H>����SBt}�S=��!5!r�{^>�g�����1�y�M�P��W�9G�l���zY3�(�W�@|���'��o���MD; �H�:��B�O�~[�B8`�CmHV��P8PU�E�>@Z[`U^��=�����2pZ�X�D��=tb�_}���ڎ-�;��jY�.\���v*iw�p8ݰD!��v4��N򼄈��� ,�B�a�MԚ��kQ
t��ˍ�VѤZ�g���>0���r�iH�9$��|]�P�`|3�tW��5��s(+�]�h�!����a@��?�(�9`$M<6WO �lD���?2�Q2wv��ɼ�&?�
1�wLw��B�Q�{�������`ןV�v��Ԍ� v�E�e�]��'݈�/�����.�ŭi�-�C3��X�~c�<2�c�b6��W0���x��	��ZV�����a덺"���� ���X�º�_��-�\:�J���t�h.c�ť��V�H�w�%Q���v�����ݪ�X��X���e���$2J[��� w��ؿ�u�i�[a4�����ܞRG�m�_d����a*jW2����ʇ��~3�3�O��;�c}���۲M��d?Ȗ7�!���W�Λ;��r ��D�{i��p[�Nr�՚ozc�k�p*��.��ֽ),��m�7r��bB7@Om:����#��	@#/~�ƾy�ч���B�6̭Sl�Wx�S!���Y$,H�!���)�X^��Em�q��郊�#�-Ӿ���5s���+��+���!�)N?v�Gw+�'�!e�m�"���Ӛ��p��ȗ?�?%F2'_ҾW{7V���ó������1���ڙ&��D_p����X��(�xp�y)�,����R$���xd����Sį~�G������÷�K`F[��N��'�c��*�*���:Y�G/�c?!J(�eIM��7�_�EFb��ڔ;���[���4�R ��`SE�bھE����u���"8������/i�v�ջYV�S�ǹ��\�s�"����#9��i?��d���b�(�r���.�Ui����a߹=@�Q�
qӿw����˂:0_�a9ß^�"���o.�L�{��ɻW��$���悼^Q� ������-�ȿl �{�㟮�����B[RL�@c�y�Q@
��&�h��U���-�J(x��z��nƅf~w֧��:��O%�0�(��[eJ=�yFs��!d���1O�uֳ�)�HE�A6��l7Y�Ȟ��c~�(f��㧉l	'Y�s7��; qt�.�k�)�Oޭ��_���� 
�=ڽ��:�U=m�b3���a������M��I�(r*��-�j�Qډ�1�8ܶ��>b�^$"4ml�#٬yU,�>JU�>#��*hҏ�
�15���/�W�ڱǴ�G����lå�߅b�9���Rd[���t b���8�ë" �o�
�$�66�g��җܜ�F��h��@��DbG�~vj:A�:��0���_���x�΋�\�Tay����
�[�K��߽�u ����y�����v֌F#�2�f�z=%���(�]�D�ދ���+|���j�*9���iƮZ�&��" �Y;�s�@v�N�Y�褟t\�-#�V�X�t����ܾezX�H�(�����~)0c��d��S�@�У�z��R@���1$���b%���