XlxV64EB    39d2     f10d3v�s�b��yŅ��$�F���N�)/"��
��{��d:F��,��|D�!�/S��7BV�/}�@�ҴK({�2��!Ę��|I�`iq�ۜᔑ>֮t�ܴ�nE�
:X;���@Ρ-��Y�:��t�ج�6�^��%�,I�V6�]��=�9�mob�Z���{�Y-'��zJ�tԺ;�3�a�fP�R������:*<�M�,zy汗�Hc9ծ1��$Js�6�C���(��x`ҿp\,	�|�_�X��@j�ʑu��i\6C��X.s{&;�ۣi1T�������.c:~ N<V� ���#[��w�Q�e�*w���a��'J�\����QT�	PhX����6&���j�1S���T*U�>�V;��\������R3����Ȗd�j�jUE׺=�^�̇��W�u�0K�Ѝ���E!4=�uf��>{�'\y��έB���O��&AFX�d����A-�B}4�'��q���o������ �Ʉ�ZsmO�"����{\0���M$����E�����2#v��\�f��`ĜJg���/��B�o�'C+xnd`{e�����|�>��La���^iC�px*��w�r�q;]���}j��q`O ����@��d�di9�>,d/���y�MƴGˉ��ɩ+���UC�~X��\(��tU�F ��
кC�OY8q������I�W�a6	�l.eE)F/���[�����������3�5�^��+ޗ���V�A�����D5J
ceQ��"�f����ư�����?�KI�Wfg�׍�i�P�Q�͎��ڟIKj?������P��Å(��J����+�q����I�l��o̶*�탵��4�2QU�Ĩ��/�~ʎOJ  }{��_@y�DBG:���5��_ݒ�QOW�>)�L�����/���a�� ,8PCV�Z��/Y6ϲ �W��ւ���CE�Kw�!B�5Ѝ<�.�a����h5��(��F��ߗ�/-a�e�����D���/c�#���C�2��V}2\�y�XYE!��cm�a�'y��J�ۜ9Dp�X`�3�Pz���~�?�aGH���L ����ّCG:{���),��۬ l�h��r�To�l+b�;�������i��RI�27 ��������:�69�S��O[e�!W�q�=�ڞog�*�Q��}�s9pА}�����f:Y~dHK�]��{�tn�`W�]j�d�ه�+o:p��}G��� t��DX���-rW�3y�[���-Cz<��T<�;�_}%���	<0�j��2�#��0{�/�R��N�0nu$H�?5)��{5���Trpv�Ze�ક����HWU��z�P~��V�z�XBd��c�~T���'\_��0�!d�}x��C_�2L�M��RB�}V��a�r8A���3���n� ����#���������&��'#���N���X?~?���ۍ`3�t�Y�ļ���Lm��}%(�1�-���Y��)"Z����a�ȃ�C��}�gZLu�e�3��д[��k����lT �8DV]�p*M'ne���ey�ӓSH��~4$����^AW�T;��y�T-7�={(.��#m�/e/�[�-��E��pkF�bL��f�s�zkSew5KH��鏅-��EG��8 �
]~�"l���8'�,^�1��e#�g�����ψ�>��^��6"��,v>��O����p��|}��0'!@[�(��a@U�~���-@7�x:Q�;Z"�D�b�l1|u�릆���?N3�e�#m���t
���͔sh����k8=����Q�JY�|E@�-�(ge��̦3���W"���3ڀ�t�fɠ?U����0�8�6T=��ȯ6:���YP���P|�sӥ��@Y<�ES�u��D�e�=cuF���@��[�%D� \RG���(�t�W:�r
I+�E* u�h;>#�ЄkG�иx�ҖZm�ӹ5L��'bd$QH�NX=��w�-I�h��n�Vr�F�=��=��8���,�j���}���6^���7Æ��<lU:me���݅vk���|�H��Nԏ��b!cr,]���v�VX����9��2�=���6o��K��$s�Г͓R��*�]�&r?P�W�Ʉ�a��Hߌ�t�s�L�m�LRc]�!S��ۘz�*���������i�	��5��K�'|߲�i�D��/n?$汅N���f��l�av�3��" e`T-5���l&]��VG�=;�r�����g����`A�|t{��\�!�ˉ�����SP����ƺ�	f�bK$���o�ߣ�L\��89��ɒ��<e�"��+cM�r��=z�wɘ`���<�TA<��HqUtL���Y����4�ˉv3����K'v�3��3<�$:M?e����i���)|w�����+g&`A���L����vMބ�O�{��0�0_Z5l&�~�U�� �6���:��2rZM��#�9��_� A%���o�k	1y��S9�f������c�k�z)�/=��_��wv$+������<3�����?[f~^�i�k��[5��e_CM�CxK���4����4��_71EL$e��5�{���]���s�>+]��#��d!��Ӝa��p��F �J�JBPa32���s:��Rt���*P I�,ul�dQnNXjnV�Z1J91n䙕ʏ��҆|� rz)���@܀��z���n��+82^ע��� �K����J�ʫ���m1�fw�a�c����j�#�*�:�י�9U�߮Ǥ��w$Y�}����ii5^�^��a�{��=XCL9g3�z U��U�r�e�7�9�P��2�Y(��џ.��AIp *�ȓ����YU��G%Z�����m P�W����r�Q�͎�?ڻN#���Lzm�������}Œ��L�����b����_�O�ŕ㙚<D�+��} U7�����v�xQS����}Q���4������=?���M��z4fql���<����VpL3~p��^J7� �>G�������A��8� #�n_��*-<W��s��� -}Q1aއ�e��E��JDQ x67yQ����.W�]�)���|qy[�V�ל�%n�1͌ۆ���;�M�5CS�|ȺP�Z�#�뢻�⹍'��{5�+�1s�h~U.�`+wVw�WI]I0l3��0"�yP��|�+��V�e��0C�B.�M"������XWԊ3�>���������!L�T�C���&��Mh�L.�p�]=�V�ĕ,��&���A0�~w����dDm�Z]���
�����*Z��Bz4�ƾx�-��xR��M�W3�w�<C��c	 0���}�;� zs�ڀN��"�J�b��6��6�,j&���Rl��}j˝����uPλ�;������Vpd�(�@xԟ$*{y��sV�aJ�	���T���f����0orވ)�>�����QK�=T�����ZŰ2�C]/~O���u��G���J�d��譹|#�6"��c��� �G���g!�T	���RŊ�a���">��L�/���S���h���'>�cUߚ�"�h!zع�������a�·L2�"s�����Pm$?KCC�'ڮ��6�AՔ�7Z�<Yf`��,̉���)�7�6X�������/�Z��Z�e�/v�Fq���y�m>�+s>����?{�<��8�'�r�Gz� ,]���*�qW ��4�Mc�Q�{<W+�h��`jI6���G���ӻ��kC����(&�ʘz4�s ᓅ�R