XlxV64EB    5767    1410�f�r5�>C���m\�>f݋�� ������ѶK�J��h���&6�����J�J���J�	t��^��K>u\݋��".���&O?��M�MRY��������D ��7n�@M��Ӭ���B�޺�|D�7�亍9�H�xb�$�V�|X�y� i����C���3����av�MR��>�y�,ܧ9m�������4#���-�$�ěGg1�bN�ѷ%�_..�#��T%E��#��1���1[2�m��E\"N@Z���ٍ%���J����[�@ʍd�@E�a��K��6A����ܣ8qgs�ܛ·[��D�=�S��v8��	5V��ܞ���u3V���GʼDt�b7����'i$�~�0&Q9�$9�U25�*�bt�G�j(��<��4j�n��9��-�[�4�!�sh��պ��m"�RrD`ݶ]un���K��D��	�r��� ����[�������.6>>E}�L�W$9����a�>Xbל�i�Jb���m�<�4�D9Ԝ�����&��\E+0��3Ne���zeo���H$�D7Zre��O,�mm�b8n;���-��*�([O}:�7���v�^��kȓJ~�r�߻o�<Z4�ho����4�˘A�"P��!���p��5���pu���?mO��mɷT��}"!�o�o�h�Kz�}�D�h�ϒ���1�`6"�H��k�Q`���,0*1"�b@��B�T7�~�_p����U5������T�� c��}�8�i�Fڦ�(�ض���K�)�h�t��D�H�f��s'z�[����G���nt+o:\Z�ͣ����c��aZ<�Ϙ�' Z}沄�n���R>!�`즇�ņ��'�o~�5L<�%����F�A-}�wgt���݄��u�)Wg�)W\,�-��8����&�)J#.��Ό樮������[��[�iS)�+�����.8�Ҷ9�YE�Px�AmU�'�$���.���dd�bi�AQ�0�8���� l����d�}�']�D�eE����]w��� H��_�뉉О��)>B>��le��+ƭ�Ό�JQn��*�N�<�%K�^�k2љ̵�l���S����K����t���]o%Xy���崍�_<���� �~��>������=կ�}$����ki^P�ٰ�:�{�`"�$M��B�4ts�]��6_N�����%�h I$G� n���*2��%�̴����7֨�C�)� �Ύ�X��������Ʊ ��,��\0����Z���O>CeՓ�*�(����FQ�A=�`��Q �|&}Km���4O�Y�s񕰽�����|~ޗrǜ�'���s��4�$8�\��Vm�U�� 3�!q���4��o�	`����n~��}K,�a��<diY��f���~^��'��5�1h����g^�m�����{�"�#�N Z�;*Vؗ�|Y|01�~���B�6�k��b��\����w��Gp9 ��lZ�]M��z���aL�tZ��z����F�P��g�?%rD�4z�������P��U͓�SO�J~C�T�pJ^���D`�+C�6$� ��2G��d�����z���1��΄Aĥh�?�OY��v$�:��������8�k��D������qyQRD9A~�ᝣ��8R��V+�)C��ǹ����M�*+X�K��w�8�t�=���7-�d-�L���W��������[�����M�yg�����t��<է�-���:��:HM��
����B1'�TV�������Z�9��MwPY`!ڰQ�l^F"��,,�2�@7n��D�����H��e�_�{�
T��L�	��)c�u7���K4z���NJk��&���<P归=,q����M��"fq�k$3>���6����^�gj��2��n���&��s� ������,�g�l��V$۹n�F�@ߛd�}��ZA
;�	�ү�&N����H�6 Fp��7Uq��)���d�0s���M%8��Y͍A.D�����~�S�W|�
qm�K��Rs�=(}�"��7Q[{Zd}Jj�o��f�A���2�m�#}S�]��EhB����ZQ�]-��i�]����R��g<���L퇿71��T+�ZEdށAm����Е�-��W8w�L�C�~�� �V��s{�$$KI���B 1� �*�����4P�?��j�n�߉�i2���
,�S%fU-u�8-J̔��������.����ۺ��K�	��*�S*ٵ���9%.��[�^�@�$9�#^�m���lq���8�b�G��s)e�7�r�[_�d��_�) -�N�DcHyO�3���o�h&�dq��{��်� ��DB�	4=���j&	�t�pc��]sza&*�M]p����|R��S5`k`�K�f��"U$Fޒa��0u}|5�^c[K3�>���$|}\}T���-��T�oՓ*2��j�x��)j @<������������IƯ�v�na9�o�@2�-b� O�=Jp�����-��X��at�r5g��wR��g�xbe��na�O�:Rřl�%p�m��S��3;㠍.C��Ӎ~]�1���zQ�i�m��Ԧ/�������M��{����S�;Y{��U;� �e����L�
X�e���xh��P��l3,�Z,[8��5J��I��9�s��ͻn~xc@�~��w<S���{��~���b�o;� �0g��BƳ����!�t�9:�V�9/"�7D��I,���g��l�G6�Te������>�K~�/�(Lόwʪ,�QPr/fO���cy���7l�L��KB�C	nX�2�����K#`\}v]F�Ǻ��f��Oh.3
�����2?C.���-i����|�Tr�v�_BʚG��2g&�x+8�b����2'8A�e���"���W�SZ��:��k[9#f9!��+ZS*��S�U������U�mA�&��t����C�[Od��e�����p%�9L^�]���K>�p�p�xS�s^2ޱ�D|Ro7�L�lIR]\���;���SB��9�m���4�r!�O4�!�a*5�[e��0B2�����޶��������ߓ	��QJ�������v�:,� EX��~q6%!Z�6��a��5��@��S��*o��77My\L4h�[����n)��i�f�k�n�q��ۛ>����ֳ�ٓ��.#�*;c��k<��ZOl���Eu��!V�K��F����
��C��jF�e+����r�[Akmխ�� �!&>�A�1���]`Z�P�~��̧��6o�f���a��Kͼ.Y��h�c�of;<@#�wZ�1��=�����SJ���^��|��ٝ�kl3��[J�K;�5����zʯN�$���p�9����j�2���I{:�Y9�CZi.ӿ�CU�@	��$��׀�SXZڲ,�K�2��T`��8Z�k���j��o��<	��5�����ќ�i6�]��QoL2G�Q�X��N ��K�0�Y��os�Gr+&H�t'��v��M"�����@� ��C��3#\�}��E���j������*�%�֢���9������b��j�7�kdrdd���d����aNDո��;T�� �~2�<�A��a5��f{x�L:���?B������������#F
%^����Q��u��W�>ڼ�.QKҰ�ĝrG�g�"ĭ���}�3��|�Y_��k��_(hO;G�.�<�!�����ȝ�Y6 '�i$�/���s��gR���6}���9�b1�
7'ʭ����h{��%��d�e�4��{�ښ��a
�2�v�âCo|ʟ�*�9=d�dؘ��@m�=Z�4VI~mC����X!�m���Q���iT�&NqWbu�L�� ����kEוٶ8U��쵭����J�&�2Fe�n�Aw�BhL1~;��G7�F�ꂺύ0���͍��L�Eg>�z�n���38� v�n�������O��ENef�\��H.��r�:?���5����G��n)���Nh�f��A+QU��j[w0J��һn���]/R^�B��m�4@���fz�#!�e|Ԁ��.6�rO��R.TY8}�B�[t7�E<�EI١��U��dtm��9�E�C�C��)C�8��8i;j���h�����8�)3ˉ�rSXG҆2������\��{����W��_*��"3�ڦ�w��]*M��0o����0�aSݧH���s^_���wl��*@P�	,(�-�K�H�.�]�,-���^f]VK��'��&��`6�������ҍ�D"7�$E��/IC�w�
�l e��ݞ��:�
��U���R"͢N<ٺ��R�ݤ�pD(�/��[ǯ��7�՝��m��B��I����QIG�� g�e$q܈�����&�+��O�`3��D�Ѭ�(��#�3,8yt�<��� #rW��'�q!(�ȳ�7����d ���C!��yR�Ɠa���>~��`2?]�%D�o8���B��8�����k�l���ZY�ޚ�S��x}�t�6���	�4� bQ.N�-)���-p.���0g�����:�r��2��ci7P�}�7k�4�42�l\�(�5L���p�<rM(ߥ��Z]�5��*G7�B��3�Ɩ���ر�ⷌ��d}� �or/����p�X-��EG�*g��b�����Ă��{+�nٯK4(l���?BF3S�����?+�Y�F�&�>�n�4y7�`~+D^A�,}�
��kp2;w��������3�jj �o��f���u���ݐ(��-ة�麰�#�}2���_���
���2��	�byG�|��,���A/[�&0v�Ze���Q_�imٹ#���9@�V��kM�|��tb��o�E7��!;I �jSJ�H$b�o.���5W��#�����bf�����R�Ō������&?S`;���-u���A���*[���*�E˩&_�e��a�\d�V����jF���4��Z����`�7��Y+?�����|��z�R��^>��k�19��