XlxV64EB    fa00    2d40�S�#T�|7v���V��2�gw���o��2k��S
GCv'(�FM�#b�N���l��s
�p�����&�cv���I�h���gB&5�wF��tն�zFǞ8�uZ�>Q�r0��G͗��0�����<�ݩ:�����%��i�~�ے0���"���.�K��]D/nL�:f����O;֦�-�o������%{ �jbI�b�����C��3����~�c��Xv7���m)xN<K������.��Q0I���"B����s�lzd9k�1�:$��Z$�Ya��O�l��o�{�꒡�H�j^����~`߃�rn�"d�;B�
��=�o8j��>0Elb���1d�ߗ�,���S��.%,ӣx��1�X����!��o��ŀT^���oL�����}K���]^�X��g��(K�PP�d��L�<��jA�L�6E�O8�d尓\�����{�Ǳ�	)+@@0t��9 �}S�q�[S�C|�^3�1�-��P ��,�:	��k�e��M�3P��x_9�*�(w	�Ǵ���F}%H�%m9�,P���V�u�i	]-Q�� �!��*5��X��~�Q<ac���Z�Ԩsx�u =&b�v3�B�J�="k�N����{�Y|�[�9��4j�������Hz J�2su����b�HD�W�<RP1k^脰`SƑ����Ӳd4I��,&���g�ٹ��`��>-�8��)[��"�K^��Rb�+��l��k=)#)B�τ�S%�&f��4�������)

���@��.�i�<3J��Hɗ��Mnt6��Tk��)=���　T �K���q,b�Y���M ұ�H�F�J��HD��Y-\�G�	vGb�J�U�2�m�l�&����SCUα��P%��h��9�Ʃ��m�|�<`�s�,�g�B^ ����43]�(����Γgn/�	W_�I~b��c?�]��,� X����ٲb[�{�!D�� ]�5��M�����u+�(���1�؋,:�1�Ǘ[�M͖-&�k��[�ו}|ײ����;ȑ���r��4������������4�Ƙ㴚��{���?��f`�7!-�^�.L�2�H`��ߺ����&Ǽv�D�m���Fob�N	Af9Sel�=�W�,��ωFw&�CD�o�Я�	�Z8�������sAF��C�}j��%��� �Ҽw!�v|u+���.b��'��_�p�S�G\�oVL�)W�~ޥ<2�1�%�X�[��y�ɵK����5�7���4���!�s���_0oL��5.ˣ�+Ҕ��:��Bc�bƽTCa�5լ�
rgx������-wT6�`G�|?�|�"�,g��ުE����
�<��6����C9B��Hd�����/).�ⓕ}@K&+�1W��K����A����H���e�SS�~�XS�R��Ņ��}�*G�n�����+[����lb�B�׏r#ô�S?E�ļ��'�X�oQ�-�03�d�,
*��+�pd�A�N�Qũp����8����f�f����`���(�b��{�_%��4
Nn��v*4P5�@\q��W|��UG�	����_\Er���䛃}ZҨ�$�J���$X��qo
�PW�dR�1/��r�Gt����ǘ~�����l���P���d�衜Ꮊ)��u��W
����'�v�m�p�b$�����4(��gU­MU��J Wxn,D1``�Z�OW����2�ߗRM�9+,�_���@�J+��#��7� �=�!m�z�j'���賊���aA�Ҩ��wK��Pda3�k#'zk݃[������-�f5��JQhb^�I-��WM�+؊[p��Cc�)����d������6�k��b�<����u9���F��[3��eo.�ą��Du�q��AP�����gU���%�*��pd�b�Y�Wl$�m8!P.|x���ϾRi�if����Em��Վ�� /?��YK�[�l��Eϛ�L9��Q;���z��.W�V�Yӏ�5���n�K犸���W����@qW��3�򀾨���/c�%R�;ŷ$<d�g��}�t�8-�_���盁��S��h�[��C�ɲ Ůǖ�4�oFs��*�-�����% �@�ԩ��-���Gs�(iBy�8 �B9Rw��#�c�O߹�ˀ܃��?�.����5�H��/�l�m����%<�^������}k1ʗU�-��ál�+a�b]��6�d\�=:I靦���wn�"��q���K7.�d{/\d�\eJd^���0>��;^� �Q����ͬu�B�s�6�B�x��,��X�w�WT�͒�k��jb\/O�뺧G���P��F�M=�/C?%�y�)b�n��Bh���q|$}�0��	]@̂�Z�K��&U?���g�U�O���W�:V���� M�5M肆��x�o�{����5�ڏߣ������\ؑF��HHr`����A���&�[��1���9)�����[) %�fѰ�n�����?�4�\�O�=U��Q�����"�N�w"0͂}��XGZ����_1,U�f�>�[����r��Ⱦ�����h�{U�ԅ�4ʕ2��ADp4�쮀�o��⃼Bqk�D3��:7�=��W[<�/�ݮ��Q��1�����s�QS��P��S-�&��ѴJ��:(� �=9�&�f�"��/I���r�}�w�ʐ3+S���J���E�|����'tP���:
�j��~6S��}�����QޜHf���`��$�������K)��k7Ҫ�L@�,*V�쵀���p�xRc��F��s&_ ��jT������K��rv���K�A����FG7&)��.ԃ`�uƲ�=翨J�x�e�[5M�l16#���U�OZ<c-��
Q��}�����$Kq!��r���A��ӎ\&{�m�t�u���<$`k\��W�k9 �%��$�O���M͂r���L?��A���l�9���f;so��>l�G��g/�{㲬�"!�L����)g\��D���k�<�L���Ħf)�e�������/�Q7�Q�]�(�i���2,MR
Tq9{X�!�� �4�ս��bDq�"QΞ0����o�Y�J
��v���h�HY�=e��GP��+1N�K� 21ׇ<��%��e�[�y���~��%���Ʈ�D��h<��(>�N+��f\�h#�!��$:wtCU�*;7���7%����q�(�U��U�e�=�G_CЯnqIq�"��2��'VP������&���a4/�S5w��]6�ATҒP~�>U�yx�b��c�]�dv��"Y��baWD�~��˥ �b�ߐ��P� �{k�E�b�9���]5��o�;kk]��-��8�Ϛ��t�wa�F6��*��������tP�K��t�g�B&�"tv�\����GߎiF������ݻtW@���Ϡ��H����6^��iJFU�(~�P�Me;IR!�Ԕ��Ҳō���$���mZ�Q�E�GJ�K��)�*����-sÖC|�������/����mȝfD������j[OO�:��P^3x�e-(j�+_}�Z���*�H�������Ǖ$4>��Ύ��{2xӺ��O����>����mr��{lD�����K�Qas���
u���\3�G��E���|?d'埔��2bq�n��s��4�G~	���#�V�T��/{�/6��:��|��my���x1����]���D�}[����^��&��FDͽ��Qt���DJ�TZ3V��zh~9�e������n7��->%&����D=KP3��S�o��?�#��1S�Ͻ���~��n�-�ĸ���{�57��7t�&�(G>_��x��x�-����Oh9���ڑ�E�uA��u]�D �:ݣ�y����oYt��E���Ѓ�G&9����5	�ITH1x>b ���W+����b�inp��~uOꭙ5S'3���H=�p�J<�m��a�T�qU�V���aG��$0�s.�dq"��Z!F�Ҕ�Dń;��6�?D�_���T���c�M�_u�c(������-�+�.��p�J"�c�|%��9���'{�:	��>�Bq����	jƲ�7J(N�_M�a!�ai�N�DP�L�.��Ct�X!h
��8�x�ryVu��6z8���-O�GLS�t��Oo�7�LVח�s������9��H�bI��0~�|��Pa�!�p��/ӕ��ؒp��䉜¤��L�LÀ� �Qz��{�Ҩcg�a(g�G���{��KV�Z @a����L�
XDz� dy׍g�Q*�R�_�{8�8������K��is���7z���f�����#���+7�!���X 9^�׆�-����inz�	��wɘ���P.�\��<�CK�~5C%=�Ŧ���_���][r��o���y�j���g� U�5�<7F�?�S#�N�*B�xX������@�l�����zi�����@uI=�5{eB2~0B�M=��h���Sx�P�?�-U���x��Ě�]I���V�è9kD�R�6!2��n7ʤ�RSKWTW���*�o���4V�j
ኅ��d����-�W�S����Jpć�+4��#@�TQ�F��uj�f3�1��7a�l�
A
��g&:m�ƍ�u?��@La�QE��ྸ��"�I���%�qZ�VE7�`]���i�1��d<M�X���6>>�ᵁbx`�etg���n�)��X!����W���{<��C�v+��d��I��;��1�ҕF뫟�$ޟ2:�S	��i�;���W�5N�������6�˶�lpF�/e���ￃ6��)_E�Le�v&O�`�0�B-c Tݳ�ꪻ���r��=O�]MYi�Я���c-I:ze�V�@^��Z[D���5k�Ѣ�6���@����y%Md���3΅(Q4ݔn Ͳ.̐lT>��#��W�@���xm�"D�d�;�I���/!��T#&c����*q ����>9cr!ƕ���V㜣$�Q��<�c�Y��)�9�UV(���iB��	Ϊz;TOw@睅�.��Q��I�С�S�I
���D����>'S@�����|lA�6,��88�0�xZ��nNb�#Ϋ�k�e�&�X����#�?���skolZ��~�-�lg7N��yo��Srqa�栠p�Im(��Q��r��I���[�ffhy����5/0������.}Ǚ�b���&.'����e������=멑�<(����HHu74���Ij燬-5n���p�������'���L�&y�����x+��iN9��8��JY���,�`�J/�iE uh���}��A�'����Dg��nZ���@�o��o1MX<��-g1�1���#�}���,��2L�}��;s�A����-�~^��g|�������K�3�^#���_��|����7�T��Mп�T�3ID�Vu�I����9��I��1IŦ�\��&9Bş���d
MQ�+Xh3�_�����4�i+i��n˱Z��ƺ���Q�%�X"J����_a5��\�u�:��^q?a�UVt�T�XZ��7!s��p��0�܁Y��-{$T�8ӭ�KżF!�r�أY�lH�v�u���)����Zo�9�!�H�w��y�u��x��@'���]���׋�8f6{Нb1��.��]�x6ҳ�^{�6=a}'�F}=C=�B��,�uKٕvS&�Ku����3u�Fj� ��m.2a�Jm{s̾L�o �N��+�|��p���+|���1����O?�5��"�;=���'.��{	^XA@��ִ\^�}
�ts�:�G�~+R$�]�(�<5������E����cā�<j苭��+��_��$�3��d�UaR��7m��2s{���`@�M�d�g����t��p�ɠ9�3�E�j�]s��ͽ�x6���p�w1˂��Jҩ����(���-�a����dn4�c�f��N����,�];�>@���Q�У���Ez� 7a"��/k+��{U�Č�S\*�(�Ҭ���a)���!��H�sK�nH��ʾzO�E+_������f{�ww��h�D���}�O'B�
�	�y5FyH`f�Mg�]v���d��_��0���`^��c6��+��\BYS
����n�ǭo��˭��3N	G�8�fC�g���)Ôo����P�'�5�w���gn��@(�5&_j?��̹b�&Z k�u�ۂ�N�����)�LM�\��W&괩fȷ���!�D�g�z�xD!�S;��i�I�I���j4����%�r����~��t��U��\rpO��9�ɤ��
D9�m������� MI���2?���z-?�,���t�y�� \����}�-s��u�?>�ݪH��PcȖ-��럐VKV����4�v���S�8�;DDA���6ϕ�}�@��Mx�����3\fIP1x^l��nl�a��k��
0g(��MGt���s���I�4�,���l۴��%��/��`����U�L�<{d��@_�Ԋϝ¡��������G�H�g$�+��6��Z��G�ݧ���'�GRA�B�J?�R; \�է^��Տ#$������yW��6n"�%��{1?�Z�v6��#
\�#E�_+K$�Agz-�MlF�y�q�� R͎(���S�<���Qf^cj`�����.\��B�k�̻��(#ocĜ�KQ��Էr���C�`�p��,vz�Ƿk�*��6��W����8wp�ք��P�T*(��&�*}�"��D�C��O$� 3�����nUbi@a��C�v�:��T���Oa�����	��,�8��>%��>��o�RQT���{dd��\��
�E�y�ӓ)�2m�5�#��|���b<s�$n�� �FR;U���3�[z�N���jip���A*��w���6{���C�X�Pk�#���6��zN�M����W�ڛ�\�*�����W�+[�gtQ#N�
Q�	�	�9T}WR��C�c�է͕)J����n8�z��,��7����ǽU�9�b�/�+�XY�G4R�]�M���VÏ`�pӤQ�>t��D����^ۡgh�)��@��HՐy�`C�>kNc�~�0�Ls픳d��ce5�;�*F�I�l}5,I�	nJ#�>�3�Z�n�k�ӵ���`^$�O�������m>��$����@b)�
�]�A��&����Z���%��_v2hg�j
>�ş�^"�0���["eK~s���F��8��t`!�hЙ�u��w�ؤ�����Ǣ��X!*	O%	;��P�lV��7�2uAX�#3��K
���xq���-] �5�J8٩�	*:��Tg�P�1���?����+"P#��c�3MqJ�(��1�3�h7����7�̑�^�@�m}f>��wS��Q�dC�MI�H_mܦ�f\�S�M\���tϮq��]:3�Ha�5Q u��8(U��o�qO��u�D�=NS�E�'��uJI��o�5��8�r�m<ر1� ���3Ms�;���4��p��`���M"���ag�:�Ř�)
ak�ȅ�jYU&�B��lʹv��̫�3�$�d���]�΁-��� �F4�]�b՟��u=�]T ��̖{v�Z	n@�P��|b���ͺ9�ȧ�9WK���]�.�A�T�֯AB�����2�����w�����Q�;K�Ѷh$��z��O�]\k�/�ЬV��~��^��"�1FtQ��h&)�3�XU�7^�k��)gU���X&�?�U�7�[��5��k_�t�k�P��!�?��Y���yˮ�󴏚q~IB\�p"��S�e�-�W��M�$K-�ȟ(L�	���n�c{����p�`��W��]��!�ݺƳ4������A�\&:Ϊ�3|�)�n����Jc��ײm�{;yc����;ߍ�+X@���)�\;��dԘ�;��Z���c8�%n�1�EZ��w�ecb�5��@�&��W���vtع�<��~.�F�6��4�oM3kڼ�����ۼn��u���B�Ŗ�jq������Ue�ʀ!��U:�`Loj����0Hj$�k��|"ދ"���ob�}�ؒ�߾`HsG��,�#A���ksFS����7B�k)`�����0B���|�@N�O��u��^�4��Dl����B4��H����T;���\w��*��<�b��o���4A�z�8�_5��^���"�إ]��''�O;�WWV��հ >�Q��T ��=V?W��y�h������l"�J�Ta�K�����ٯR�@황�M�r6Ă]��ڜ�|�t��F��#��ow�o�ג��]G�\V��:\��sϴ�l[�RDhqֽ2�d���7��4��W�<lRj&En`��p�leCP��?ٽ�N�L�[�M��{qYv^�ѱ!�����՚R��]�2S����^��<Ix���i��.g��v��59>{m�ǃ�\�O|L�y����pL(�i���%|��PI���@CT�}��;�ئ	>�:{΄#q1�5�~�uO�?[h��*����W&Я�/`��A��+-�з��p�<��{�� 5�r����垍����CmJ�;�Ϣ�L�C���\�!�������x6qJ�;7BE��Tc@�]�>q�;�Bt��U�r"p��uB���� �9�Eu�j���l�x��'Y�W�uB2��[8��pQ>�����%�)��0�c3w�ml����$t-�ipk�o�dG�����K��]v,'����	.��Z(�0�}��PK�3~)
F��F��$90�\�z�+����Lt��\C��[�<���:s�`G�>f2�X
�;����;~8q��=b%�[�~��ǱN�>I$`�b/N�yOKT���lP`z�Q�h*�fN�@���)��d����'-M��և��ݓ��{�rʱD��+�-!BA��a��6��}eGn���i������4���>CC�����"������%�$��3�������)k��z�m�e�I�� ~�k�t��L%���_b>��� ��R*\g
�-��Txic=�V���d��غh��W�����χ��e���'��4�A�p�y�q3(_F�0��w�[�����s3 �;x�2x����ѧ�\��,@�q<uL���
�κ+��7��lHW���p�z� 6(��X���zP2��j!��BӥNS*���V�,Ki�&��g�S�������p�m��OU�Gѭo�����a�~�����ͷ\�����O�C��$m%�ɨ�B_�ߟ�8+�w�3�����.������G��'0�R���p]�0*�k�)kTᤳ!?TU�>Z}�+���N���X�E�eΐ�r[�`m��������3������
bD��)��YA#��X%`��;g����	=E�Q�Rp��:!��.��QL�����LC�[��嘚��y��k>\��}r�������j���>�Fo�N�g�\{� ���nDۂq|���w�A%�&x�[��1m�/FH��_�v␥�{�x�8Q��ae}$ K��uF�ob���=H�y��,�
��W-8���夡��XАn�����!��J�0��E���G�����2]���B��`�44u�m�lܹ$�����}�H��h��ѧ�o�1sr�\s�F(0��/�/��y��{�ǣq�xԮ�f	gF��}��B1�z}UJv�/t���RҢ(>_�3`�!����Hj�8[��A� Ֆ�=Ŀ�R�5Օ��]e(�_l;!���]��<��#�}��E�p=(��-�V�m�C�<K�|\"��:;l|h�]z�D9MA���t������f���}ꍹg(�8ʸhHo��7�d�V��ں� ���߸�T�#�:֔7_��*���l�����<?�3c�2򼴁���3�#l0�dŞ3Xm�G\l�Xqes3;_Y�_���$�*G7����:�m-���W�,'~^b��9�HF�C��N�}�k=~�DS������-e,wԢ�?�ka@����bo��i�p�Í41�XJ��p���%q;��f�<S����_|	mƚܾ�p���Z���b�IR�bE�gި�>����+g�a Ƹ��f�E�["��c�7�HՃ�h��g�@�n<���Yړ�=?��rj�
UA����fuG��L|1�e �@Å{"^x����F-���:�ھp�1�����5a��=S�ۉ� ��PJ&N��߶����{����x`&�����s�kJ�	�Y�Aw��_�;����r�cf�ph-�(�=��Z�d,���|&�vq���$Z<ʃ�#��V�gG\+8����fv���6l粸u�z�
L0��(��=�'^�~�,�=4+(��~~�]Z@�v|� &��2���}g���<z��������C·%#��G�e���K�N[�X��۫�#���w�����I�3��l�V������<�.{D.�!}6T�a�Љ5�=m餃�G'���5u�꾂�(t��y���}6�;�h��LQ�ЈI�-l �Q��+��Tj��*�|�P."���,�p<�P֥F\%4xLT�AqA����>�$$T�#Bsυ������M��#�M�t���w���h�Coqo�G� �0',�
n��y��˞6v����5���M�)��t��m�����PD>6"�j@��ckQ
}�D7����%��%r��KAaZQ 	</+����X����Yj�.s���d��
����n��gZǅ?g2�����s�U�&"�H�jTν�nx�K�#u���)�ą���������8�(����z���6S�T���Tp?<���MZ��
���6��o`�k�p|���t�~��Z쏤^]A<e|6���.�~��+q}�c8B�6
��7��8m��wE��v�%�l��������W�	j�.Ԍ{{s�":��t*��Ts\l��*�|Ni��j"�a�0�d�����9��,ΘDg]N�����9~���#a�sQub"h����Y�Co�/ķ.:�Rx#0�\�ˇm�`&���*�V��;>�A�����ӿ8�[���w9y�l��ә�.p�)z�@}{G���ɢ���R����{�F]w�ݠ�8 P���N5R����%Ȃ(&^m��:�H�VHT�T���]
153^W1[�$�Cr=�_�Sۙ��;$���|<���è��JMŝ\c���[k*��ϗ��7nA�Х�YD�
Q�tz�Ӷ��x�z�P�5�z��������V�~]�(����0�o����SՐ>��zȫF�@ޟ��;�������rZgb�k����+$����[���p������o���ѓ�\bF�d���Ո�XlxV64EB    fa00    27309
�ڮK-\$���{�tI\\\a���!�.�'[�_�*�ifU�����c�}n�[�A(?Ƞ�f�4|"p���G!�R� r@�Fa%Ē�B��u�~�1�H�OuNqϓ:�-�
4%����]Fb.A\��4G|h��q����+�Z����ݭ�Q����!��x���z��Fx�K4P���L��ⶢPDYuѵ�yR����E�΍K"<�`e ԓ��D)c�%+��U%���J�����c��q�-k㶘����ɾ"E��(��t%�a���`2��+k����>y�2jU6|�Pǃ�'��&ˊ�1l���:�ۨo�Ǧ���) �|tYr�mn���b�����9pR��$�]P�|�z����ѱ��
���f�;���`9���>�m�&o�� .RL4���Ss)M�Ŏ��V�+��0��UD=KdE�s��+���`��'Y~5�� /�ܶѷا�`ą\��&�ލ�D�'�e|�.+�Gm7�Q'f�|� ؖY�,)���L5���d!!f|���p���PQ�E8�|Un�o�H�w�In$Z���~:�/��4qB�6�M��:(�u�?[6�>\�f��,0U~�5���_��չ�'��V/*��㎣]�[��e��R�I��&�����/�����"Z�0s��|�F�H�����E���������<}U]�v�$�	�Hg�$@ �H��pݴm�Y��j\c����68J���m�ݸ�վ��k�:�&w�暖Rs����tc
Sw��Vu)�ح{͵='״?�Q�TH�p��`�u�4�7�y�V=H�v45��%���:��ˋ��
�� n�z?�e���, ����`�Gs�J���6^�w��vFBJJc�}H))vZw�}�m@-9j�>��۵s�M�(rL��N� ��% ��@y��醌��XO)�����B֗u�\�`��Ɍ�]��7����i�,�R�s>�i@��E���6B���ȇ4Q�S���KX�}P��쬆<� �C
OM�@w����[���)��rN�9N�a��H��� ��@����yWGP���0	O��)���=LXz6�!�����ͨ�κ�蠬�a�r��y<�݁�݂��0�~H�>7 }#�u��E�{)���MDl�@�k~!��_%�Q�A/5d�C�q}�evn�3j �HfR�C�@
��5��� Rդ:��T�R�	�+)�,���y�b��$��o���Q=k�#r�MҠ��4��`����(N- �f^�Tц�GV_`��S�5c*vi5��t�蚫6]�IUU[�Ts]5D�
G�M�(b@�Deq�nV����
!�b9@�)��T�H����`���}#��oD�,�t_Ub��k14����'+��.������Y��#Ƃ,2�#{��v�,Ըo&9F��ʚ djf@٫,�c7��I�Hu{��]����PG�d�9:���5������8�p3�
$.w=�%f������^� �$ueEeju��܇�E=�3��#+���E%��[y��TE�KKw�)��g�6�o�M�q&F~`���"�1�l�IB1B��~)�f�07�����F>g�~�9�֔�?��9U�<��0`O��;#�0�6�&yu~5T�~x���Y�	��*�֥��2�:ߵKJ��X��*�O��ͱs�n��.2}�.�b���� N"o�]��/��Wg���SGU�����H}���3� K��BR��������+��,�$=�<j����*_@��ٳ��1�{�&8/u,~<#�|Zl> ���z O$�7]$ǝ���b�[�?�C���k`��������˯����`���iq|��ό��є/B�~)�<�.�CcD��fXx�}'7��y��k�$��0o���5Ʋ��vm��R<���2������{�A��͉4"Lȝ~���6��Zv�)�#(��t��YF����4�����+�Z�M�7I%���I�I�TĤi3秊�N�ȹ��cSsYX�.����4x��ǒ(r�]�MˈEs$�!���F���E���hC��*���s� �2�:�w��bq��Pb���0�㳄Vܡ��WR]�EΞ�,E-��{��ϩ��w��}��i���N~���څS����p5*vH?i(X"����xb���V<'���/֍|�h�x(����+�߷7��� �[K������Y��D��@g�z `\9���B8(�DrH��oB8�&�z�9���-ƨJ,.��d[�ɉ�p��;��H	��Ń�owZ~.��V�����~ ���U�_\��B��-�/,8��5m�n��;Фp-۲�EͲDڥT���=ӌa��d9��-��O��*�
�����\���p0���~��I��ϥ
˰H
b�+�� �q;�/�MI#���Uv��ݥ�J��+)�K�;n+I8�E>��&P�7מV��d�>8�Ղ�}�T"���.��3��]�5����j��7��0r�]���I��`N���r(��D�L^�>��j�X�����B��7�?(^S���dx����*��􍳒<���\��G�:�ɕ���0]E�ҍ���W�~
p�D���L%��<�;`��t�&c�����f�;�h�q��p��2��ߞ�Dh|�����pz�h�7د��=����ʵ0c4�#JS�d�&D���=b��,�6�_c������=��Z0��b������#g�"�ۂ#�*g#�?|��)~'��ęG��u�1V��x���j&�3�=���i�l<Xs�w��d�6h�#�]Q��Ĺ\��nLؐY }	Q�	ax��X	�=i
]� �z�g��]J���tt��1�dr!�~4Э��'0_�7�Y�#z+�3�t+%���|�#T`�r��]~/���z.@�T;]Ol}l6�cpO��.�@�J�Z=�:&�ֶ��j)���3͒�P},��E������V�L�BeD�H��*a>W�e�c��]	��Pr��*^����t�H'�R!f�ٰ���������d}X�Eo���$5��0��_L^4�A�� �	�i�|o�]d_�ס�=�+�f��%��e�B��#n��R�F	�D�2�UQ��|7� �Ծ
z�#a�F���{�ܻW q�)��
 ���	z�At�@���Kq��������'%�7��B8=�/�W�fu��U�%EǸW)\qƃ2l��xO���-/i_�A�� s��R� �GI�n��������|)�eVՀ�3����C�������H!	�j�m���8�IM��%�9u��/T��e�c�	F�ެ�F�hM�Uߤ
u�6�7$ߢO���G~�V0q R��W��\G?S���e���;~U39M�t�)�����L5r����}J.��Q}w��>/F}c��V����@Ѹp�|!�|�2�)$7La�T[��:U��UY�Ykk��B!���We5�, 6"4�=��I�m<D���?
��p��S���N�FJ��n� �]��:+��q�@��C�}���B��u<�OvH�3�i�+<B�o;�@3��VO2дf�A?�+���"�_v�%Q��&
c˱���Hi�[XIޭ��=�KMwFS �)˕1,�| �`EX����3�3�ԉX-�4��&J�r����b��Nb ���?,{���Sa��D��~��m_�U��<�%j��W��&a�>��F�l���d��YJ�l�H�MI���#�Ev��$���S��*��ۊIDs'Mn|۬�I]j.��w�����bI�+|w�m��m1.[O����iPi���5?�yn*�Q�����+'�W�*v�=3�X�&jKr�`��BQ�"r5�[:��Y�{��������Ȝ�J���z#��n���O�I��o~yt��/�7���W��RQ�]�'�b�����z�#�5�?�*:�f�ƚq��fQ�.��w����#�sZd0�����a���B�u�A2�6MwYcm@�~2�Pxƌ�>���-Nj�D�n��VW���Zi������n}��NȜ��c�U�����S}T�V��Z��%�፦Q��d��lJB�1'0A)�pѥ��y�	+�16N�m��?[�~��y����_��Y��-b�����;����"�B$il���~���O���H|�'��	�Ky�iy�W&T�p"v��/b�D�Pe.n�H��X�@���f�����g�R�n,��(b9�4P�aC/p߈��lkh�ɍ��3�xD<��3i���������V�e z��Z�E��w0CV��f���9��k�+,��2��O}sVmV�{h�t�ec����'��nj�C+�	�!�@O8�7	p�8�yƹ;��tSA8ʳ �v1�Ќ)R��-�oXu=a�yqktb�>��g ے4v�O�sph���4���`V�_L2Ǘ/+�m��p���9YkƚM%�[�U��f=pm�K�,ڭ�ϲ�Wg��.U�6�����}�Q�UȰo�%/����{��I�v����׊�Ŀ�l���;!�)�w��U���ob���/p�Q
Qۘ����>1���l:�>T��A�d��
k��N��QB��\�z����� ��T1:�w;6��.�Bx}@�_�E�3c���Yy�Ӭ������Xp�(��3�}�Rų�U�L�p�H累�%�B��L���
 �uy���߽62�i1�(D��PV5�\v�#��cfÛs��Zc��[��mn��}��gxQC6A9���s�LV5�-� Z���&u[!@�� ���,�cz�;QKڕ��d�Ԃ,�"����}u�|4(�ɞ���f-���$P�J_�:wb>�Z����X��J��<Oz��	]�J�U��4[ޭ�y�G�l�є�]HȲ�[ƽ̩��� ���$��+w(�:yE��x?X��q�q0����*�?�>Ru���e4c�<�@(����{K���i�'�q�M��+��5\��7���� I�i滋����T�jAK�,a�DQM�K3`(�h%,���K�V�Al����[m���b|�S#с��6��ID+��1^�yz�P���!�c�V�*�V�����P��5?��U�ٌR�|��U���kn莗�����\U�x�aDXK���4:���gk�Ð��H+��z�F���K��J��آ��{�s1�!h��,�o"/�׉�M�	��?^6��uE(��pl{oӼi�Fl�k�!6p=.ԑ��M۴�!]uc���m]wE�B�� �J{c|#���؏w�$������I��w�ۺe'�~R����d�5]��/��p{���t3l�w���8��E�a�c9��XO��1�ۻOS����L�8;|ՇrD,�D��p�ʗ�|�z b���eN���"�@�VBS��	#�aA��X��	g$8rI�j/ȋ�y7P�W���Ցq�]4�L�!��"B��ia�ĩT	Hy�rRm�Y*�=;7�y�|�$�v��P��|{<5T�-���QZ7�C�g/�������[&�%�\�Aº�Bz����n�UYY\�s*�rrE��s�K�A�*=e�).X����$�=r�����h��~���0�i��b~�O��\
�kz:K�V?w�ƣw��=|V&c{j	�Ў,.����-ӄ��vn�JD���U��0P�)z�<�B�.�9K��G�0۬���wr�`?��o:Ij\��֊�ݫ$YA�#">�M�E\nWG��\�5������W��'w�	�s����m�^a�D�&`���!�j�i�]���u>��ƥ6��ѷj3�����:�>�{B�}��dR�Q���}��4e���C�x��Wj7@��:L�a͑����0'}w '��=g��w�D��Y�J�G�^��L���"8]��#�̺���~Ҏ��ls��w�某�2[�_/�jE�y"6�z��a�/~Q�%2*�	ŵ'�^�n�Y���T�}�Zm`�w��f�	�Z��4}D�X��ϲ�T +�=���7��!�>y�I��'��k��M�[��ՉG5t����.����Į-���-��1�
�~���w��,�z�ےBQr�T�Y|'�]��;��,���'ރc�-��B:�L)����Y��)��K���![��3s���XJt#j*�n>��2sYA����/�]ˈ3�2@u��j��)=˱~�=�gK��0��?8�k���5���n#=¨S*��x����f,=d�����(�&��4���N�b�#T�p*ຣQ��@�����uDΣ�Nx��lڞ+���}���F�h������O�����M$�f��n�^�����g	�S�$�ȇ�����sQ���~h������!2�*�(]v_@�-��zL�a�<�Ռ��\��2L�l0.�>~͉��E�(+�c����a�A h!$���َ� �4���ʥ�|�b����'�m�طv�5�l����)#9�� z�R��\{<������N,�t:�޸�J��~+]��'G��J�fn$đ��b�EX��Z�5�K*�i����7�Q��&�1s X~����&?�t�S/Z��M�IOG��Ꝿ�/p떭�9�ܾ�f�~b�=�?b��w�<W�߽�;�;�F����h;Q�Ą�Y�}����(!zD�9��ƴv�D»�n���ػ׀����c,n+���'(�[3E�A��$�6�k��Av	�-�=�
�#��'�l��H��m�Vuhƀ�\/pN��v���;�B��g͒g�|���٭u���Vq=�2_[�, �^Ǎ;ԑ��oSDj��lER4B��,¥������g1.f�<�~�&��yg얆k%����=�QV��-��Z���P�԰����C����rٯ1G`nIx�R���LXȌP'W4e� ����6���2x�!��c;Q[x@�YIH���UPXN��*�yK��+� �~¹�W"}u��RQ��&��ư����i�29q/s�_���]�JY��C���SF�I�a7���0Jú,L𱼘�X.x!�2���a�azi�	%N�|u��r�dW��+�s�D
�2�_�_�瞫uO���;i�6wşU�h¸M�I�x�i�@���:�����fX�.gu��Θ���}��&��aV�4���z�wq��[��_�VN�	*0~��1	i�-=�U������B>�������; ��1�;(�FHjc<E��-bY��6;v���}C�]Mk�M�C���{�m wc������#� �4_/Y��+x��l�C�,�Wy�N#+�t!@6�^���Г�~<��ߙ��-�����HP�<��A�'�8f���{��GGnzN����B:u����"������+�	mW�>L:r�	���AfoM�I�G��T�4����[P�fk ������������b����|��,���pn���`!��oX:	�v�)�Ԡ7N���z��EO�C�g��J����E�����[s���й���Ey�����[������|����b1��ǭ�0Z���)�����Hi%t���1�	���%�Nw/�=l�HP~e*����J�~n!�+������մ�S�]�}B��1��`r��G0����&�	XTT/�ߖѥ�m��Bϳ\��$��g|������,���Y�ߴ�/.�A��j7qЕ-���uZ7�-�0����)Y�@��τ��.��8N�f�{�C�@��Ye�RI����=��H��HK�k߉;��1���Y(�q/����R�|�e2�c�;�AqMO�O
��"8��,S�\���0�������O���M�O@�Ӓ���	�0\���QR�ɵ���6H,O�3�*�f��>����հN�2J� ���k<�*D�t5��T�H����ዡ���BX5{p���a�ں�W��4�����
+�T��ѹ��ܦ��N�g�p7��:y�;���d�jJ�L�%RJiÏ"�a�y���\qD\.�Z�mT9����;�?���h5`O+7���Zbf�@���:#hQp�_�wr�	NAҩ7\������n�|��Pb��������a���y�`��LRH�6���'��Kې6�$q�;U'(-�(j?�E��d(�B�K�L�5���*E9���ӄ<⪷�A���Z���m�3���7�q�g����
[iH�o�0gK��q�i@ɛא��w{f��,��#.(�o��#t�PS.�½��]w�T�A��?�L�2� 	�S����ࠋ,��'�U��QU��EC��hb���%���@G�p�ʲg�Ǫ*ͳ��a�y�[�Q�@�q+��S
��T_���v�C���7X*��&z�T��v�����n{}�5W� >0ʼ�pI�.D?�>/����/G)7U��R��y&��nf�\���owh�����+K��
���\�~i�E��+?�LZ���h,�(�]�W/�25SWw�k����$����e@���W�o����坽ߊ �t�
8��Z��&��ڌX.���=�/Z��}6ILp�$�<S֑|�$e�'�c?����X�`�Wġ�àQ9�����"�{����s�����6"���|	X��'���!��k'xIwS1/��S���g�z#��g�:*���\��'�;Ihg��&��,{O�a��psɤ\����0��Ҵ�8�-N|�i�_ͤr���.�\�mSt����6 �|^��o�z�w�,�>�yS��8��-�x�}o��É~��=<Ze�ߠ�z,}K��|����߽g�7�-����ⶇ� �l��������N��ÚȑK_$t�z@�(�gI�p���Iɵ�$l����O�c�J�o��b~s��i>�I�M]���ȫ�'���3���A�����c>c 0�p\ .�*��?���:z���hd���Y���cg�2딲Sv����V�Ȃ'k�}��J�ˡ
~��Hl�F���LŠ�+ՊC�����4�VwE�zM����[�9ѵ��7k�母���-����6�1H�������.kO�����V9�;����m�^�>؊U�͉CMߧjna�CZ�����k���X��J�����	�XE<�拥Ev����[#����A�a�a�瑖��:�p�j����6�Xu�o��;�=&��[BF�K����L-;���d��z���}H�d	cПƠ��4r�jd��Fz���c0��5��Ӹ5�8�)�r]� �5<V9���:.YH�)bV��eo��br)�0�I��)���ۍԕ4��qx�>�_�@�.)���~XB�iTf�a��3�6T��AK�����0�`����֢�Y�P��c�]/`ƺ��|�x��P���ڒ`\�(�҅G��-UC�`S�}����,ޑ���ěm�Z����zX��H��� qh

)�gl�U�� ��o�I��>�h�h� #A�<*��|�B(�hM:�P1� {��c���ERs�橉�,���
�������Ivf 26���d�	�^���2�d��
���ܢ�*g� �cd��elڒdd�t��.��%��A�(>6z��_NW�>��/��yӈo^x���!J�&�7DAo� Q*�:K2R)F�d�Ľ?�鷏�L��g�RP���'��]G]҄���e��h8�Y�U��У�]��
.�θ��ʒ���ooj��-�!�w�C`�r�b�`�� �:��F1�K�k��=��	ȍ Θ��2RU�u
X"���Uy�������wD��f�9�'`G4�
�U�e�	�G���c'�=\m0�gq_��!��`�>��uP|復�����j�4?�����'U��ӭ1�xL ER�Gv��B��.���i$���U����,�@j5C�Hi<$.׬s8j7�XlxV64EB    5e8d     f80��1.���c(0sq�b�pD�a
�+��|\�'�������伎D�g"֞�H$�������Q��5~�i���A�h�h񘭻iG�Z=)�I9F�j!瓛���o���$bnJ��]4eGx).w>x��	%�w�@P;@�3(�kC����E&l�M�.�n��lE��4|==���$�HF��
Й�L��b0s��+4��/��	�Ͽ�g'j����4P���l�FG�}b�����os�&1�����a�	��0���|y#�iP<\ ����5��)K'��x��@�4��ޏi�;��zj��lc��uѵ$]�� �o��8",�&�.t�&���gHV�^>�(��1،��7�y�$6��6.,}H�f��@�`�xAx���~�a���C�1�i$��p���ü��@���c��BՖ-F�+�/sӲ7a�`��~i3�����U���7_�/�]"�!���)&�Oku���Rl�!�[�x3̛i�N�gP��"����g}�ʷ^��P2 �o(�8)����MK�׸�V��\Znc�� �"y��GM��k�Ax���� �.@=�k$���)U9�1���v�}��qYْ*)�씑�7T�v���~M�d2�����z��%�y4�{���������K4#�V6�A�81�ӅCBr?O�,��W�s[��^%Jb����<�t^�#���t��ׇF�7��b�8
`�c*�0�O-�QI�W�Ҥ�x��r ��T!12�pQ$��c��cZ��P��u�s�젫:j��_m�3��V�k��s��p���s��(��?7iQ�[��D�����[�1h�⼗��7����<�^P���NF��	$�k�w� ��*��זM�hB��;]�{O��Y*Ʀ�U������i$�꜁�:���ʅ��W0�Š!C�����D��a,V�i�]�c��ȁڊ[���ל����c�#�	8�U��Z�'���*���YEh��0e�G�Q!��W�(�t��$�DJߢ�QL �W�@Mٓ~;-0ߋjՑCu�2�L���?�� |]6g�l1+Ł6����򚶦�o҈�VRV��o��F'sD�D\�Kch����]�����iO��a�I@� �o��+te�fW]�oy֩�G	)`�o���[�n��)-��ld$�[��������!�'"�x��$��sa�,��5[VA>�u�Y���bZ(m�Z0)������	OxA{��u��C�f�5��Yy޾�Ca젤oMc�}�5����i���I_���[�6�X���A�z��C|Q���ej��a�kW��\�*.%/�������fC�l�ǭ=П!@Ԏ�z����p�r�
��t�CC���\�YF	X ��@���YE�G�M�$���:=��7��P��
�Me'vt����]�j�V���
9y�+�,����-��k[$1ĩh�����ks���g��"N7|����'�:ũ�|4 ���5���1�0aO�D����L#1w�u ���g�4�ꯀ�%/��2O/�H����q�R�OMc��>=��W�=��jeQX�^�[m�M�E0����9�� ���w��J� �����niGIi��e�^O��	�3|�+C��]ӑ�����l��"��}_��~C�����C��������Y�9��:F��cf�l��#�&<�J6Z�,�#��}�FYX�?AH�p�ڲ ^����p�-�u:���*�ϩ�pkM�)�@�9|K��/Xp(T+~[�ˣ��l*����]�����`�18#��߿�֍�Bf�����G�5dB S�܍�*.w+�u��4o��I(W"w��J��n��	��������:�&,�t[ZKq�v�ѩ�/�n)�EO:G��Q��i_{t,'����c�,a�IF�BH�*3��l�52��I/U�Ȫ�Ha�S�QVM����
�Ac��(��"�K2�<���3p�C��"��*3��`�Ra�c^.�x��?@���A��}�C/z�^$��,<L�Pr�v�_����enB���B9di��Q��TK<˱vI�$�V�_���B�OpO��jV	S:�����5n�N����AOt�è���CbXX	�^����zLe�������T��?穯�aʴ����X�7��ț�cx��:��4S9^ 8����m���[ht闗B\98Y������܄��/޴�ՙ��H����N&�����x�		��y �%�d�)D��j���W���C%
��[?��*#��l��x�UB�v�M&9I��i?�m'C�)����h5;�hb�4~m[��S�v8������?�L=�l�[8њ���u#��10�ov�Z[M���-4>d1&�+��H*�T�/�\���9�@-�P� ՗:��e��q3��n*s�������퇰Ie��������f���Cz�+(^K8*�,P9�c�u�4����-�Lb�u������EJ��"�P�!!I�����Ri{�IB޽�$��9��2K� '��˗��ƀ��ږ�G��0�:�O��WY��ͪ��gi�}"�	ܼ��K�J�ʲ�k�1�Qz�{���ƃ�%l�s���8^�3旰��n2�m�KF��uvxu\��!�W]�t�L_6@��F�.���[)3�� ��{e�,��5b]�F%F@1�R޸s5�*;56��ē7��_��T����|���_�xS�a�� ����H,?wI:7u,^=mm���m05���L�V����	f�����|�!�)����p�+���`#
/s���>O+~��m��M���Vi�3�x5�#5����M�h�k��i�k�|�j��i�'ۙ/���0���-T�K�������0/K159MO %@b�"	1��4`��/�g�t�:{�Pl=��d&.EΎ)gu�=��Dַd����n�VK5:#+��0�D��|� g��5V�1/F0��0�W�Uj����������Fti�To�ȷ#N<�+x��6���<\r��l\�ʲ~$AB�����W���
mv?���?��AR�:���T��vfܙ �LI��o��A|�1�v���<]�/Gyz�c�l��_�@혩5ѥ���j���6��H��3��q��>8�
!t$\xL0Uf_�*����ކyʇ	qv������[��c��Ԓ���F��
��'���+"�f��U������G#�<DeO��?�u*t�2�T��fq��]�B�k�-`
�F/Se��D�����v��u��i[�SR�$�
+�)����m ������w�[;��m��[$��h#s�EX`;��i������;��f��x��w�5B�Qe9��wQM�`H��A�Y�	g����!��I���e]nζeaH�AVf��0�g��(����Z� -}�~c�y�@���?��]@ȤP]���r1��c���C�������.j9��(�K��5�S˅���{,��ǒ�Ϸ��t��װ����g�: �[�>Ɔ�.�����r�V��O�^���S�	-T{.(�F�o+�c�<P7�5RP��BX��x����s����B��I�9v\d������P��"����
��\�"��a�į��T�rS@��������Y�=���/�z	%�X��ĭ�WY�of�v�} ���`o��ݻ��8p�]p��K3j�qs�:���s���{�v��{�49Prxt�}?�v��\���3Mq3�}-��0x �B;�Ό�B�V�*l��{Z-���( <u���
�6���u��޲2>w��B���7rpu��[B��M�<��P�M�9�~%�����iI��ZpĬ�A��nԢ&�[�&���Q���L�AT�(��"k2�y�RW�\�=����([&�#�R�Sf��H`=�1���*G�?