XlxV64EB    346b     e50ûХ�۫J�o0>srk\�
��J5�P�|.;�bz��k��*r�QG�E�����tO�	��jB���
���T�	& ���C|�R��K�k�z�VD>7�gæTS���d%���>�e�A��6h�6��rUG�G���ƳF�0n�;�8�O���=�E�_z\��`����3��+�5>��?������i��"䑑�׫@rY�B�^nD�Ȗ�	���<8��~��7O�?�~����㸻];���5S)�E !ph�+�J�nc)'�C���8p�=-�haY%�\��jXh7b���1�W%Vˌp�*<����CO�O�b�A���t��'�R���C$9�2��+�@M1{��M�A'��ý�$��Q���$�Fn�#�ڔ,��s�)�����F�E�F$I���F��o"J M�ݙe�(9*��:Xc�H�vc1��5De����V����y*0�����>�_j"���2����+|_��ҝ����ٍM1�1*2����I��J*���w`=!R��r	B�տL��9?{BIdX��~Mm;��j���u튫�E9"��@�jM2!��z`/���ߚy1��O��r�u��z����Yv�9n@�� �o�e�����Nb�3j(%Ջ!t95�g�^�rZ���]���-8�"�������ּ&c�:Pz�V$�q�p�<P��� �Z{��K��%�������/*�fdY*OJ�a�X�%��AO�/`Hp��= �p$OXE+0�vu�}�0"�\>�Z���\y��7�T�����!�TMh~������w�/�q�6yIX`}Q�k����ձ���6��Ջ�sZڳ�pK�� ��)��K;Aߏ1/!�#dTs��[���9�Б�Oy,;o�'`�����4����S�l��a�>��C^F�'�Ǯ�FX�?r�6��b�"<��^��������3�aח��<���F,��Xr}3;�~C����\܍S��t2��]l<n27��������[� �6����eb������4c�s#�Q
���h�4��� 6�\8�m�m���"Vy5^�����D\O_�A�Ν�|@p/|�_�xW����v��tD�+@e�s ��#��W'[�D����+ݵ�QJ��|����J6=<��I7Uhu��"�ߎ��R%W�I��@yp
Sq�wزcg��B�� _�����ÁL�!͍Gb���1"�l$�u�7qm��
���̧�H���N_5�!�i�s�V�&���ű�ɯ+!���,} ��H�֭��XD��+���r�Q��gY�&����h̂��P���{I&�t'D��RK��s��^BL.R.q���U��{8I�؉^���(_��Hn�}G�be��iM *k�W}�X�1�!P����:>��Bo�9Թ;`�"E����A�XZT�fb����T�&��U�(�g �6����XD����W�-Z�!��p�'7�	�
�F[�x?�YK���Ӑ��~��ө�}&M��xx��y�'+ia�('L�5-ͯ��Vl.w�J5֚K��� ��]V�ㆢ�������6B	Jo|t=��Wf��5�a�A	�2S�s�I��!sJ�<8�����z42���*���Tv[�]t���#	P_�_�ԋ0�'f_{����G�O��S�<��� �$�.v������+]�v�Z��Tk���/�d��X_���Ԙ!�ۺ@RF�fC�}T�u#��e��1�PB�}4�B�i[��@��ʻ㖅s�M�G�h�sbV��j�g�2�ؤ^�~#Z�53��LgU�,^���d�D9h�f�`ʟHC�J_�{_�9+�߶��b9֧�P�~�|ˎ��V٫=H�Q�o1ܾL8k�e��$f�q��d�y��F���.���O(�۲	��_Ͷt-�b$�=�b�Ԥ�}�8� ��4;��Pa�ȕB�$�|�}�F��՞{��6߲��
�����R�~;S�b<�P���G��-F�p_l����Z>��16��M;�c|�ւn,�ќT�K�<�u��W��m@�8eG1�S�uck��U���_#�s��r|u���o��Bq��	p/��x�S�Z%�^5�1�M�Xm�*��������0��(G���y�-։;���s!	���"�l,�'�o�1V7׃c\�
1�ծΚ[1|}��D�#Z��&XՀ8<��IVBApE/�i̵A��'�)�q0s��
���e�s��[+��4��$��b�mpb�x�y%�ŐRқal��YB>�	����(�j�cmO&z�� �4)3���y~]4K��~Co(Q0`[\���gGX}��j9a+��\�{r��l~�Qr��a+�2�����6JK0��OR�s�h!�mV;�PL:���	�-� W���tQ��aj!E��\:�C��a��9�v$+���m�C����av~��/��h^��Yj;�e��{_~�K雘���xt�E�r�IF��rBi.�}�����
��$�؝�ZG�ۆ��M�j�89�t+G��p�P�?ok!N�"x�ֈ��p�_=�:`��J}_�����,w����lHǋU`<�J���d�gu=��H�y%7�f�;���\���AJf�v3����r>��T�_�^`��'��6I���X�Z�]U�X�}�fZi��
��N�ua���#n��(��}v�I�w�M!��Y4�|t�qaf���j��}'��
sr�h�9��m�4	���tS�/�u�Z�E	���� p�R=f<�rQ�3|B+��pl�R&	�_j�F����V���||��GXrG�������՝j�,�y�'A�u��Q��"	�	p�Zp��������/ ��_h9���%k�{lD֘�����㻤ꕉx�$y���R��NA4�	�XN��T�kM�����-q�਋�'�����Q��*햂�f�į���/�f�T���NF��~�UԌ�<��^�@-ڬXLLbd��h2�ǚ5n��3��+ר�6�Ś����N�Z���Zi��ū�.1o��v ��}�e5>OH�rh�6<��I�4�'kVpo����dJ+B?'��6w$�!���54%fKȯ{���*���_U�	B[ &]�{�Od�5�?D�n���J��V��kM �՜ }@!Z��S�Oó�sZ�L���<�K���Ds�ߋ#>� ������eG7䊽�`Bc`�t��G;�������	��*�yE�� l[�I��ɛ����M�3 �Wѡ�����z�Dm�&�|��A�Yqõ��S��R�[�NjLݽh��=sf�y���I�+���i2.j$������9;P�֜�Y�h!G���.�A��_sf�"<`�/�L)�J.|JҺ�����A5 �Z�y�-)�3�+[A���|�#��F��$����w�[|A�*z3K1�uU��K5.���[�4\��B��wӚ��`(�3ۧ}&�x��	3�\�%@2����f�$p׫�5������c��
Ņ���͐2"T�d��\2|&
I;p1%+��G�xS�` "t`O!�|��I kXG@��@&g	g����B�0F���b�6k�`oC��"-@����j��%ڮ��!v��Gt�Z�,�Mm���y�g� r