XlxV64EB    21be     a60�L����߳�A�)=����ף����`;�&,��t��f�x:�;��L�S�zH���fu(e��C��/��/8N�WD�⿽���@uɢ~c+�c�Ⲧ�7.�V@Q��|�[b�WE*n\���z�R������>�kR�*�}���05!d��8tὭ.L0��
N�jj���,��b���~�I1����)hrC_���/Zb|k�/��c�1A]]&�����:��0�FPw<�G��j���9���S���J��P�i opD���uݟ���r@���Ԯ�=�BNu��O��s�~D@�k�o����
��ɟ�:�SޮԔ���ߒ4�>�d�ʯ��\��?iI��ܚ���4y�$�b�{�+9L�@<�;�P��xW���k_�]X��9�cj<�7�)�$��&-�v1��(�a+F���*4ԡ���^鬈h�[��"����m՗��1[��$/����^�T�ԧ�_ڔ9��Wu[e��4o+sq.B��v&�\/�=�7�PӸ�b2&��"���?��h�@�u�秓��~�Rڲ&�%�)�1g��)�����Ϸ��CQԳ?���W�bG����a��UO=�D�~�����9�����)�qtI,�g���t�܇;�����S�.�m� cP��Z�
�M�'	�\�ȖoX���%�j�j�:�[���/q�ݛ�K�GK���[����X��u�7[��P�E��ʀ5a};��2_9��f�ڣ��{F��z��:���NM�W�X��
�ܬ��KU��T�=Ȗ��G���,R%������4�'^-0nP�M�� ��:X&�	�p������i8���y� AOQp�уT��s�Κdc�/GƎ��o�Pi���@��u�kRSz�v��C��S�������3�)mlL��c~��d=sS��:B!�+z�F$�g��@����zP��%���F�o�^
���bPx���fݭ�la���,��BT)�7t���<3�迈��v��gF�a���E�rYtgI�p���}v���i!r��ϛ��7��5A���(�H��Q�3Wc�0Ͽ������Ɇ��i{�r8PEU70���P�KL*S�ڗH��QhD�]9_Y�=8�s�t(�"7�7�T]'����^Q��z/�>�?�a�����CT��ZQ� Yy�1�r���*�ߘ�D�t	���S��5$�a)��}m���Y����o9��D.�Tʵ��� G.�M1:�l	zL�)�:_6��!I�o�u7�K�������`7���k��P6'�1���^Q]F�~k�dnn%?��W_*���\}x��<뜵P/��t3�;���6f�b��ɝ<Wy��5��F�7s����VT��u`�]��+6������-k_ƺh7���]K�i
\�{��.���V��u6�=�W�� �N��s���W_�G�B�Ix��#�ѡy������ �ި��d8�����p��N`4NM&-eU����bs|����o��I	�+�]�X�^CoL���s�K�N�Ĕ�0����I֦��9�4qo$�=zZ��Y�FʽDD�Fv�`��G�'���+�=�7����T6:�m�^!k�-ֆ��0w_YP��c�lr�_��RD;Q�Ď��=B���7�JT�Q�c'�,#|���6��/A��0���ȗ�kV���x��x��$xԔ� r�������;���hJ& �wwD]F��iϣl�Q�}�qOq��?4�jF�>b��f+�ʌ�\��\f�J
��/,��^��ŎB��7�������|���جx��xC�W��]�w�guA�R���kl��3��Y�V(�*�6�
���h�����P�x�)KV�yl�1m��>\�Px�;0$٬�B}W)Eu:/��MY���es�&X�*� �1��:h��s���yk�,��<�,�=���2i��N_i�a�Ja��S��Xh�~�J_0�3�����я4���W�E��r�g�|u54FO�$CR�'VJ�Zkc���Ól䩊����F�˲�ň�VhP���_>��2��(�o�����kۺY�g�Ϙ
�����m�C�����p#�8�D8h�Y�<�IN##�-NllS5�m[d�b+���H�ʚ��[ƈ�����n�j%�-��<!p��V���ե�=���#�-�&�Ӓ	"ϟ�W����\�ؙwCs���&��蜡C�$�wZyIވ�$v0U�E��Oۉ�(�5�=m	s� �`�K��.��lt��� HB��
�ؗ��n�p�vm3C��/~0��L5 �fX��WL��Gu�v��A�l� ����Z� �p�?����X-��N�;(�;C�d&\i��-��ƈ�/9��N�+l����`� �143�%`Ӕ����v�w��a�s���ӋC��A�1md�3��x��9��,���n+��(�o���澐qh�e�0zq@Ⱦ�y���9�%�Oğ�r Y_�Ƣɛ�^��}�ﲁ�"�b��1��9lcpz�X�/�5Ju��|y���[�	��[����K�#�^~M��|���kA��5�W)����i&O�7�U_��eI^ ��_��Em"O�r0��N����%d��N�)��(�d{���a� �c��=Q�����ޝ��