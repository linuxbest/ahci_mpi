XlxV64EB    a7b4    1bd0��T7ބ���8Q�;�!g�ը��g�U|`B5խ]��˧XS%�A�3)��ǠKh�jXd̽���8����cNv�`v"�W���e�98z�X�@�8��W{�$�$�*B�X�$'\��QJE����7���Xُ�m��O>�Ѕ�����8�+;�.٧,}�*Pm4Ej��J��F�z��ذg��\�^�4�HTg�qܧ�0�!H�b�P5����>Sx�{��v6t�����9P��s]��s�b�㩞|��p�j*s[��˭Rt����(�]�:-�l���6�j�%zb�zH
�Ěhj���E�9h��*g-��0��Ѩ����&J����${sfJ���2�LU�3������q0�L��̎����ŀ���	�������y�d¢���M�3�3��	�䮥H{�;_k}���'V�0�`��{[�C�5�:tE��o�kX(½�*:Sq�s��{�t8J̲�E���^���Um�D_�u��2�XL�f�˳�<��m���05���[%ȝ�t�y�� 5�,%�!D�"�2�����t_���`�69D��-��I���*_YGO
B@<����aslx0�pj�|h��[zL�
�'��.y���7�d>4�C�j��@�nnxQ�Sf�e���^��~��[������Q�ޑ5��M�J๐5�瑠��A+�^�����o��M���]&K0;���C��È[i���gM�G��ZKg��!<��'�[Y������c ��4������cg��B�����w"ԕDL�M�Y+�~/��;����V�k�h(��,�$r^��Rs��Jʽ��\lp=:�M_���_.$�����̈fO�H���Q�_<1o���5��_	Ë�e~����n��VؤO��=�@�<�=��A*�@Η/�;]u}\5�6�5�/����E�w ޤ��;��C�;N�����x���Ƣ��e��Aࣤ��a�����=�zF�������m�諍��@�pJUТ�6�-"*>�փ�ԥ�.�ot�����v���ԱI��9V\k�/l�$[8����^0Z������n����GV�\�ƺz�U �Q�Ƴt�qz��Af�%�מ������]d��]:^����X�?Y��e��F��$�S�\�+�}��MZ� 1�� wg��ƀ|o��q����ЫQ��̧��8���rjl]��u��ap&�L�Ϊ�����:�]R�"�k�y	ג4B�m�V�Jj��ƚ"r��P�m�˫�i���R�ȞPk��E9v6�Ӯpw"([�� �@�������
�}G�J�
%��A�������~B�w�:b�-a�O�8rȧ��E���n�R��.�Ԥi��\;�������H�l-��G���I����$�:�����,А��p$ˋ'����W�m�8� �|��(��~!x����+�vigE�����&�QF��N��~�ށ�����<��}:0�il3�p����>Y�V��VV���wE-1��TL�G[(�9k�Mʃ���S��#%�������B��H���6��Ѩ��RR�`z�< nOtdg�/�Xm�yw ���JJZd�6O ή���|9L�>�GL���N�ZO�wF�j*���{5*v��W�Dw=���y�BP�`׻�:�D������+��xK��/Ο�=�ЗMۂ�s{C�[�wF��Zb#73We���� �����?L�R�- ����-O[q7}�?�OL�L�f^�^��o�krMQ���N�c>���;�k�cfUQ�^���px��~�G�:�mK>+>}H��Z�	�"o�����Zr8��;OEZ��䵛�E��͙�\�ʴǏ�Sbc���9\�e:�ʐ(J��`")a���T�������7�v:�c)ϳ�9��ѯ U���M��FZ��`b3)�qߞK�ߍ�jsJ��վ�\�h�JvAb􏆚�y����}w�1�ȗ	�����a����W���@e�:Մ/�'��fOJ�C@��/�q1�4#�J8-#�[cH`҇�:����u������X�B6!F�.C/�(}�r�K!�6Z�-���)Ҙ��)�&�1�.�jC}Sd�k�z���ɸ�\�1�ލ���5��kV���V{��.z�E�s�����	'^ lO�|a�'�i�ceqAE���-s����Ѐiܬ��a_����u@�������L���z9�+;���S��w0U��S�H>i�����TJ��Q�jO�Rec(2�9�'�?l�ad���(~��(�ْ./j}����Ā�Di(I�~9X�t�� ߿8Y:��5���걞>�o�7����Ƒ�e����h������eyN·������Mŋ55����䜮�"����pU\Tm������D�3��ߪ��}�GJ����m9LJ�mLL�K���{'g����c[K vV�](����9��N��ܶx�����:��YT�.�j�����D'��h/�m�([=���@�Sg?lI�] �V+dՌ4��.	1�A���y�S�*9��d�R+8��\�+��L!��nI&�E�;����|�խҬ7�t�ȋ���4�+�Wvb5:���O��B[���#��*��X��	nfo�ɩ%�汝�kU�B��f�Bv?��~�
A��P@N8�����z�֏ϦL�Ģ<9����S���1��vx�]C��AOO'\���Ȭ��<{�_�2D���OX��g���k�	�m��pL}m�7�#k[��~2�8l�\�PnE-�  ��p`>R��Y�{�
���"���Z��s?�p��G�4��g����k��>/=׼D.	-i�z#ǜ�d��+�҇Կخ�4���uE�碬.	k�W�>����H�XK�V����#��;�k��/�[�Onb���sZ_a'3�:żmQ��D�6䶧�N��O<��1^Wf@�ui`fBiz%x����	MT����ۻ�!/v���Ho$��Cf#-�f��AF��t��(
	;H7Z���?�;�%^��Q�z��RDzCDÀ»߆f���v�:}�H�!|��_0��t*܅�S�0�I��L�k�U��ʭ��0b@=^����
�1\���q�+�����e��G�X�ѮdoS��BU3�7PD7�Z<���;b����H]���xב '�*�>-���Q�P@�|�$9��ڎߙ��O�ե��Zh�A��>I;�-\5� hؖ��܂�ݧ.M���Q?��iuI�\� ���q1?�H��K��x�V��[pr���|�����;<�	C_�V��e�w,K���!�[{�����{i7�%`Z�r�E\�"��>��˗�ZFתl�V1���� ��|>oȱ�?%Q-�R�.S��2�Jŉ&�5K-.�(��Y7F��J��@�ّ�����t�{�L�C�[eܓ�4rĸB�����k����i|wZ���?GεF=ў�%b�t �i���^�(:����ݴ�m��\�����k����h��g��Ca�̯I3���U�]�?�����8���(X	���j˦�Z��l�7��k�x��W�������(%��m�l�F�*����"��� 0�)�������M �)�#�gnc�?儥 �*w��Ra�}���H�P b���L���}���FKC<0�N9Q�$Ķ�o����H]+��� ܁���W�-?� c�6�e����:��e�Ow $�]Zΐ��c!�V�ՍOU�Nr:!;S�����ܫ��9�݅��3z�ae>��1|�Y�a"�Tu7�Z65��ǈ)]db|}�N(���i�OQF�YԻO���2 �Z��ܗ1fn�|d�XS������x�		.cnx�9]�� e�(��I�N�[K���^R� k�˖��u#�j��ۨ|L5������g��M �\w!M&��`��?e�u�0u,#�#ye�˟�P��c�R)Rj�<�� �se�+U��(t��nS8��bH�iA�d�����n�&�9�'��ǽ�$v�#��������/�ƅԪ@��͘�)�ު�u�?޸���� %�S:��Y�T#��\�m*��$����SԔ1m����S�f6R0�V�!O7��k�c~\7Я��\���E��JsO�����_Gn|��E?�����-�|�j���#�h�ބ�1��pVG�p���~3�;�8�1�;V�x�|�?���<�y��L{k�P�8�i�Ϩ����{�M��3՟WM���Ga�sLҌ��@��^��cU�Ӹԫ��)?}d�ʎ{���C�5������ɲ�!�Y�z�Crm�M����a`�^qˣ!�ೆ�\���mJ<&��oZ<pp5ǅyd���݉�(2�SآMI� �*�Ja�*��)���)'>�മP�ȶ��9xT!~�É�5|о.�)�����/��u9j|3����<�"Mm��ua���_բ44R�J,P��J���s�Wat�~!�4�I�"��<T���T�5�McʿU0U6�D;7'��皞˽���E���AϜ;��Ƿ���4�;��?"���P�g���������Gn}L��Ը_�ȠfY��Y,�J,�%6��*���W:L�W���b�dK옥���Z��Yv؏E�$�ڧՏ���!/뷳%���ؐ���o�&�dc���i��U���p�Y!���]Ad��'������8D��TQ�i:0�4��	���P�:i(�ܚy�];�W�/K)�J�+������ΖL�e�3Yfu�9�IE��N��?�m����4��ؽy�Il8�	`�TF~M節SZnVLFH�����D�|�jɂ��ԡFs���C�pl�q���S�vg+X����[#�|j0 O"�p@��ъ�g����m�OM0���e7�[�m%6E\�R���8��x-�+l.��g�����OO�Q�Q���lr��#���sxף���sl�u��}����5$��N��p�G��*-����b��XFn����"*�KI�TWF	�8�@�u!g����8�ʥ$AU��l~�;/��^��s Ѥە��'�������&㻈����e͊g���G�9��z?ElL�U��=/�A����_�p�c���~����߯�S{'�VW�/��l�G�=�\ܞ�]����� ���1t�`G��ëG���� �s�-�5�~��A	�EHK��\��}�āqu�|`�:^�B��f7�C���魬q�pE*jW�*������ 9i���a�����V5��`N@h�Q,����;�k�����7�_" 5��MN�`�D�V�\�zc 0A~�2f�	�y\�e�P
����~.w�����Y~�[�t��ZM��2#���0.Jٙ��-n��q��(�e�=l1Ӆ�� ��Jp��-P;���io�N:�eHM��Qne:��T�U�c:%}���hq���G�K8#J��9��X���Ef
�͍�}�]���;������:ct��m\���$�v�#�o��	FuH"�i����ɩ�ٰ�&aI�ѧ}��<":'bʚ��P��x��LX�7*�`�Xנ5�	�j�Qb��T����U��u�X�[�#zW�-k�1�?��~ϟ�2�43�6n��F�`�;���j�z�
o ��t_�F�$E�]��t� ֶ\3��{�G����0 ��m���� �֦zn�����~��/�^���
)����7(�J] ��9h�:���Q���� ՕN�Ġ�p�v��Sۈ~�}j����=��������n�N$EjoHz�E��T=� �ߔ.R�TEv�*!&��K���������Q��d���\;�����j���a�H!� ȹ�k�u�/V�Y��h"*hU|�5H�ֿw��(g�����]͂�kx*Q�4Z#�n����E��#�|4l���du�l�"A�S�2�DBd},Ȟ!z9����H��S71ʂt}�Z�}��5��-����r��zH�#@%��y�_	B�?��9!*�\�W�%��_d2�ED�o�WŌ(eSqp�	���-�r	���+����q�q}E��t0��O�-9�[��af�X.4#���zÆ�MF�����u�w���3���&y=�Z�)�<Yx{�S^he�kHZ�>5H6�AOlR�+�k�V�~�pvn~ۚ��:R��V�7?([n�"������IĦAj]y��F!��X'�7��o�󺴛�:�/7)/6�)'��d�Y�J*��6ku������-=�~B��"1��.��#*ns���$�?�
�˳��'i����"��:<N�\�oɸ3w�-}�L����l��b��2*�:?_I-��M�mD��`m�_Kf���e~7:��=/
Kq��o!Ц�7U�l���¢�5U;^n��Z�_i��;�q�6P�Fz��nͺ�����(솨�+wEI*Z�,� 	5�-�j�g'fo�	D�[��ۛ�g�٢���[��6������g�@>�4�{>ʐ�*'�۩�c-���3��C�z��x�I!���B��3g�-��˩��4��Z��o��L%��SG�����!=o���g�$A�dn���R�/������(ꔍ���}�g���p_@5#��,�#��y� �
�`�+��l�5Q�ٹLM�`��X7�n��o���
����a���R���;�c�8bű�'�.}dUۍ�g�.<,�F�Y���~:���z�����<�u����.#]��XK�-�� t쾏�m��j�iDهz�:�\��aKT�='���\�8���}~]� ��zx��=_��m��v�F��I�&��j�~A뚘M�Y�]��/���_�Bs@؀۠����I��$5�[*��;ѕ�i����Ң�Q�)�@M������9�MK�ד� �H�ھy��Wm�z\.�o	Kwvq�Q�9����ʧ���-��d�������D柜��cث�i	���������rCL챏M��l���Ju�k�Λ�LÁ������i8���}+�W�B�E:�q.��k�2�2�p�?